CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
32 89 1032 744
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
32 89 1032 744
144179218 272
0
6 Title:
5 Name:
0
0
0
8
9 Resistor~
219 255 103 0 2 5
0 4 3
0
0 0 608 90
2 1k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8953 0 0
0
0
9 Resistor~
219 255 202 0 2 5
0 5 4
0
0 0 608 90
2 1k
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4441 0 0
0
0
9 Resistor~
219 255 310 0 3 5
0 2 5 -1
0
0 0 608 90
2 1k
8 0 22 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3618 0 0
0
0
9 Resistor~
219 624 121 0 3 5
0 2 3 -1
0
0 0 608 90
2 1k
8 0 22 8
5 Load1
10 -14 45 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6153 0 0
0
0
9 Resistor~
219 489 310 0 3 5
0 2 3 -1
0
0 0 608 90
2 1k
8 0 22 8
5 Load2
8 -11 43 -3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5394 0 0
0
0
9 Resistor~
219 381 310 0 3 5
0 2 4 -1
0
0 0 608 90
2 1k
8 0 22 8
5 Load3
7 -10 42 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7734 0 0
0
0
9 V Source~
197 57 166 0 2 5
0 3 2
0
0 0 16992 0
3 10V
13 0 34 8
2 Vs
16 -10 30 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
9914 0 0
0
0
7 Ground~
168 57 472 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3747 0 0
0
0
11
2 0 0 0 0 16 0 5 0 0 9 3
489 292
489 157
255 157
2 0 0 0 0 16 0 6 0 0 8 3
381 292
381 262
255 262
1 0 2 0 0 16 0 3 0 0 6 2
255 328
255 446
1 0 2 0 0 16 0 5 0 0 6 2
489 328
489 446
1 0 2 0 0 16 0 6 0 0 6 4
381 328
381 339
382 339
382 446
1 1 2 0 0 16 0 8 4 0 0 4
57 466
57 446
624 446
624 139
2 1 2 0 0 16 0 7 8 0 0 2
57 187
57 466
2 1 5 0 0 16 0 3 2 0 0 2
255 292
255 220
2 1 4 0 0 16 0 2 1 0 0 2
255 184
255 121
2 0 3 0 0 16 0 1 0 0 11 2
255 85
255 38
2 1 3 0 0 16 0 4 7 0 0 5
624 103
624 38
56 38
56 145
57 145
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
184 7 240 31
194 15 242 31
6 Node A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
181 143 237 167
191 151 239 167
6 Node B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
185 248 241 272
195 256 243 272
6 Node C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
8 149 40 173
18 157 42 173
3 24V
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
192 444 248 468
202 452 250 468
6 Node D
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
1245414 1210432 100 100 0 0
0 0 0 0
1 58 139 113
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 0.5 5
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
