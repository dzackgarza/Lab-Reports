CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
110 160 30 200 9
32 88 1248 733
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
32 88 1248 733
144179218 256
0
6 Title:
5 Name:
0
0
0
7
7 Ground~
168 297 351 0 1 3
0 0
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8953 0 0
0
0
12 SPST Switch~
165 504 333 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 4208 0
0
2 S2
-7 -18 7 -10
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
4441 0 0
0
0
12 SPST Switch~
165 504 243 0 1 11
0 0
0
0 0 4144 0
0
2 S1
-7 -18 7 -10
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
3618 0 0
0
0
6 Diode~
219 468 288 0 1 5
0 0
0
0 0 1360 90
4 Vout
14 0 42 8
2 D1
22 -10 36 -2
9 Channel 2
9 12 72 20
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
6153 0 0
0
0
10 Capacitor~
219 432 243 0 1 5
0 0
0
0 0 848 0
5 0.1uF
-17 -18 18 -10
2 C1
-7 -29 7 -21
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5394 0 0
0
0
9 Resistor~
219 378 243 0 1 5
0 0
0
0 0 880 0
3 10k
-10 -14 11 -6
2 R3
-7 -29 7 -21
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7734 0 0
0
0
4 VCO~
221 324 288 0 5 9
0 0 0 0 0 1
0
0 0 1616 0
7 SINEVCO
34 -2 83 6
3 Vs3
33 -2 54 6
9 Channel 1
32 11 95 19
0
29 %D %%vd(%1,%2) %%vd(%3,%4) %M
0
14 alias:ASINEVCO
0
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 0 0 0 0
1 V
9914 0 0
0
0
9
2 0 0 0 0 0 0 4 0 0 2 2
468 278
468 243
2 2 0 0 0 0 0 5 3 0 0 2
441 243
487 243
1 2 0 0 0 0 0 1 7 0 0 2
297 345
297 318
1 0 0 0 0 16 0 4 0 0 6 2
468 298
468 333
4 0 0 0 0 0 0 7 0 0 6 2
333 318
333 333
2 2 0 0 0 0 0 2 7 0 0 3
487 333
297 333
297 318
2 1 0 0 0 0 0 6 5 0 0 2
396 243
423 243
1 0 0 0 0 0 0 7 0 0 9 3
297 264
297 243
333 243
3 1 0 0 0 0 0 7 6 0 0 3
333 264
333 243
360 243
2
13 7 0 0 0 0 0 0 0 0 0 0 54
11 Ubuntu Mono
0 0 0 1
507 310 521 327
510 312 517 325
1 -
13 7 0 0 0 0 0 0 0 0 0 0 54
11 Ubuntu Mono
0 0 0 1
506 248 520 265
509 250 516 263
1 +
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 100 100 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12401 0
0 0.3 0.5
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
