CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
20 0 30 100 9
34 93 1332 746
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
34 93 1332 746
177209362 0
0
6 Title:
5 Name:
0
0
0
30
9 Resistor~
219 816 354 0 1 5
0 0
0
0 0 864 90
2 1k
8 0 22 8
2 R9
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8953 0 0
0
0
12 Hex Display~
7 863 179 0 16 19
10 0 0 0 0 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
4441 0 0
0
0
9 Data Seq~
170 1060 90 0 17 18
0 0 0 0 0 0 0 0 0 0
0 1 1 1 1 1 0 33
0
0 0 4704 0
6 DIGSRC
-21 -44 21 -36
3 DS1
-11 -44 10 -36
0
0
49 %D [%9i %10i][%1o %2o %3o %4o %5o %6o %7o %8o] %M
0
11 type:source
5 SIP10
21

0 1 2 3 4 5 6 7 8 9
10 1 2 3 4 5 6 7 8 9
10 0
65 0 0 0 0 0 0 0
2 DS
3618 0 0
0
0
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
12 SPDT Switch~
164 186 134 0 3 11
0 10 3 10
0
0 0 4720 0
0
2 S8
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
6153 0 0
0
0
12 SPDT Switch~
164 188 164 0 3 11
0 10 3 10
0
0 0 4720 0
0
2 S7
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
5394 0 0
0
0
12 SPDT Switch~
164 187 195 0 3 11
0 10 3 10
0
0 0 4720 0
0
2 S6
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
7734 0 0
0
0
12 SPDT Switch~
164 184 222 0 3 11
0 10 3 10
0
0 0 4720 0
0
2 S5
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
9914 0 0
0
0
12 SPDT Switch~
164 189 252 0 3 11
0 10 3 10
0
0 0 4720 0
0
2 S4
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
3747 0 0
0
0
12 SPDT Switch~
164 189 281 0 3 11
0 10 3 10
0
0 0 4720 0
0
2 S3
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
3549 0 0
0
0
12 SPDT Switch~
164 182 306 0 3 11
0 10 3 10
0
0 0 4720 0
0
2 S2
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
7931 0 0
0
0
12 SPDT Switch~
164 181 335 0 3 11
0 10 3 10
0
0 0 4720 0
0
2 S1
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
9325 0 0
0
0
4 LED~
171 407 364 0 2 2
10 10 18
0
0 0 880 0
4 LED1
17 0 45 8
2 D8
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
8903 0 0
0
0
4 LED~
171 450 342 0 2 2
10 10 25
0
0 0 880 0
4 LED1
17 0 45 8
2 D7
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3834 0 0
0
0
4 LED~
171 500 315 0 2 2
10 10 19
0
0 0 880 0
4 LED1
17 0 45 8
2 D6
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3363 0 0
0
0
4 LED~
171 544 289 0 2 2
10 10 20
0
0 0 880 0
4 LED1
17 0 45 8
2 D5
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
7668 0 0
0
0
4 LED~
171 590 367 0 2 2
10 10 21
0
0 0 880 0
4 LED1
17 0 45 8
2 D4
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
4718 0 0
0
0
4 LED~
171 619 340 0 2 2
10 10 22
0
0 0 880 0
4 LED1
17 0 45 8
2 D3
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3874 0 0
0
0
4 LED~
171 650 317 0 2 2
10 10 23
0
0 0 880 0
4 LED1
17 0 45 8
2 D2
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
6671 0 0
0
0
4 LED~
171 678 295 0 2 2
10 10 24
0
0 0 880 0
4 LED1
17 0 45 8
2 D1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3789 0 0
0
0
7 Ground~
168 101 423 0 1 3
0 10
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4871 0 0
0
0
9 V Source~
197 70 370 0 2 5
0 3 10
0
0 0 17264 0
2 5V
16 0 30 8
3 Vs1
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
3750 0 0
0
0
6 74LS83
105 739 231 0 14 29
0 10 10 10 10 10 10 10 10 10
17 14 15 16 13
0
0 0 13040 0
7 74LS83A
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
8778 0 0
0
0
9 Resistor~
219 678 394 0 3 5
0 10 24 -1
0
0 0 880 90
3 300
7 0 28 8
2 R8
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
538 0 0
0
0
9 Resistor~
219 650 396 0 3 5
0 10 23 -1
0
0 0 880 90
3 300
7 0 28 8
2 R7
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6843 0 0
0
0
9 Resistor~
219 620 394 0 3 5
0 10 22 -1
0
0 0 880 90
3 300
7 0 28 8
2 R6
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3136 0 0
0
0
9 Resistor~
219 590 399 0 3 5
0 10 21 -1
0
0 0 880 90
3 300
7 0 28 8
2 R5
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5950 0 0
0
0
9 Resistor~
219 544 389 0 3 5
0 10 20 -1
0
0 0 880 90
3 300
7 0 28 8
2 R4
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5670 0 0
0
0
9 Resistor~
219 500 395 0 3 5
0 10 19 -1
0
0 0 880 90
3 300
7 0 28 8
2 R3
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6828 0 0
0
0
9 Resistor~
219 448 394 0 3 5
0 10 25 -1
0
0 0 880 90
3 300
7 0 28 8
2 R2
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6735 0 0
0
0
9 Resistor~
219 407 397 0 3 5
0 10 18 -1
0
0 0 880 90
3 300
7 0 28 8
2 R1
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8365 0 0
0
0
66
9 0 0 0 0 0 0 22 0 0 2 2
707 276
707 417
1 0 0 0 0 0 0 1 0 0 46 3
816 372
816 417
650 417
14 0 0 0 0 0 0 22 0 0 40 2
771 276
816 276
0 0 0 0 0 0 0 0 0 5 10 2
816 240
816 249
0 0 0 0 0 0 0 0 0 6 9 2
816 230
816 240
0 0 0 0 0 0 0 0 0 7 8 2
816 222
816 231
4 10 0 0 0 0 0 2 22 0 0 3
854 203
854 222
771 222
11 3 0 0 0 0 0 22 2 0 0 3
771 231
860 231
860 203
2 12 0 0 0 0 0 2 22 0 0 3
866 203
866 240
771 240
13 1 0 0 0 0 0 22 2 0 0 3
771 249
872 249
872 203
3 0 10 0 0 4096 2 11 0 0 18 2
164 339
127 339
3 0 10 0 0 4096 2 10 0 0 18 2
165 310
127 310
3 0 10 0 0 4096 2 9 0 0 18 2
172 285
127 285
3 0 10 0 0 0 2 8 0 0 18 2
172 256
127 256
3 0 10 0 0 0 2 7 0 0 18 2
167 226
127 226
3 0 10 0 0 0 2 6 0 0 18 2
170 199
127 199
3 0 10 0 0 0 2 5 0 0 18 2
171 168
127 168
3 0 10 0 0 8192 2 4 0 0 44 3
169 138
127 138
127 415
2 0 3 0 0 4096 0 11 0 0 26 2
164 331
70 331
2 0 3 0 0 4096 0 10 0 0 26 2
165 302
70 302
2 0 3 0 0 4096 0 9 0 0 26 2
172 277
70 277
2 0 3 0 0 0 0 8 0 0 26 2
172 248
70 248
2 0 3 0 0 0 0 7 0 0 26 2
167 218
70 218
2 0 3 0 0 0 0 6 0 0 26 2
170 191
70 191
2 0 3 0 0 0 0 5 0 0 26 2
171 160
70 160
2 1 3 0 0 8320 0 4 21 0 0 3
169 130
70 130
70 349
1 0 10 0 0 4096 4 4 0 0 33 2
203 134
203 135
1 0 10 0 0 0 5 5 0 0 37 2
205 164
205 164
1 0 10 0 0 0 6 6 0 0 36 2
204 195
204 195
1 0 10 0 0 0 7 8 0 0 32 2
206 252
206 252
1 0 10 0 0 0 8 9 0 0 65 2
206 281
206 281
0 5 10 0 0 12416 7 0 22 0 0 4
202 252
286 252
286 231
707 231
0 1 10 0 0 4224 4 0 19 0 0 3
196 135
678 135
678 285
1 7 10 0 0 16512 9 10 22 0 0 5
199 306
199 307
355 307
355 249
707 249
0 1 10 0 0 12288 0 0 11 50 0 4
407 258
385 258
385 335
198 335
0 0 10 0 0 8320 6 0 0 60 0 3
620 213
620 195
198 195
0 0 10 0 0 8320 5 0 0 59 0 3
651 204
651 164
200 164
0 1 10 0 0 4096 11 0 7 61 0 2
590 222
201 222
1 0 10 0 0 0 4 22 0 0 33 2
707 195
678 195
0 2 10 0 0 0 2 0 1 4 0 2
816 248
816 336
0 1 10 0 0 0 2 0 26 48 0 3
544 419
544 417
590 417
0 1 10 0 0 0 2 0 28 43 0 3
449 415
449 413
500 413
1 0 10 0 0 0 2 30 0 0 49 2
407 415
449 415
1 1 10 0 0 8320 2 20 30 0 0 3
101 417
101 415
407 415
2 1 10 0 0 0 2 21 20 0 0 3
70 391
70 417
101 417
1 0 10 0 0 0 2 24 0 0 47 3
650 414
650 417
620 417
1 1 10 0 0 0 2 25 26 0 0 3
620 412
620 417
590 417
1 1 10 0 0 0 2 28 27 0 0 4
500 413
500 419
544 419
544 407
1 0 10 0 0 0 2 29 0 0 0 3
448 412
449 412
449 419
1 8 10 0 0 8320 0 12 22 0 0 3
407 354
407 258
707 258
2 2 18 0 0 4224 0 12 30 0 0 2
407 374
407 379
2 2 19 0 0 4224 0 14 28 0 0 2
500 325
500 377
2 2 20 0 0 4224 0 15 27 0 0 2
544 299
544 371
2 2 21 0 0 4224 0 16 26 0 0 2
590 377
590 381
2 2 22 0 0 8320 0 17 25 0 0 3
619 350
620 350
620 376
2 2 23 0 0 4224 0 18 24 0 0 2
650 327
650 378
2 2 24 0 0 4224 0 19 23 0 0 2
678 305
678 376
2 2 25 0 0 8320 0 13 29 0 0 4
450 352
449 352
449 376
448 376
2 1 10 0 0 0 5 22 18 0 0 3
707 204
650 204
650 307
3 1 10 0 0 0 6 22 17 0 0 4
707 213
620 213
620 330
619 330
0 1 10 0 0 0 11 0 16 62 0 2
590 222
590 357
4 0 10 0 0 4224 11 22 0 0 0 2
707 222
249 222
0 1 10 0 0 0 7 0 15 32 0 2
544 231
544 279
0 1 10 0 0 4096 8 0 14 65 0 2
500 240
500 305
6 0 10 0 0 4224 8 22 0 0 0 4
707 240
319 240
319 281
203 281
0 1 10 0 0 0 9 0 13 34 0 3
449 249
449 332
450 332
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
1312660 1210432 100 100 0 0
0 0 0 0
1 66 162 136
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12401 0
4 2 2
1
791 284
0 11 0 0 2	0 67 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
