CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
20 40 30 100 9
0 71 1366 768
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1366 768
177209362 0
0
6 Title:
5 Name:
0
0
0
39
7 Ground~
168 145 354 0 1 3
0 37
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8953 0 0
0
0
6 74LS83
105 808 177 0 14 29
0 37 37 37 37 18 17 16 15 37
6 7 8 10 29
0
0 0 13040 0
7 74LS83A
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
4441 0 0
0
0
6 74LS83
105 816 452 0 14 29
0 37 37 37 37 26 25 24 23 29
3 4 5 9 28
0
0 0 13040 0
7 74LS83A
-24 -60 25 -52
2 U3
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
3618 0 0
0
0
12 SPDT Switch~
164 288 344 0 3 11
0 37 30 37
0
0 0 5488 0
3 ADD
-11 12 10 20
2 SS
-7 -25 7 -17
8 SUBTRACT
-25 -19 31 -11
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 -1 0
1 S
6153 0 0
0
0
9 2-In XOR~
219 501 214 0 3 22
0 37 37 26
0
0 0 624 0
4 4070
-14 -24 14 -16
3 U4D
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 4 2 0
1 U
5394 0 0
0
0
9 2-In XOR~
219 499 268 0 3 22
0 37 37 25
0
0 0 624 0
4 4070
-14 -24 14 -16
3 U4C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 3 2 0
1 U
7734 0 0
0
0
9 2-In XOR~
219 503 319 0 3 22
0 37 37 24
0
0 0 624 0
4 4070
-14 -24 14 -16
3 U4B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 2 2 0
1 U
9914 0 0
0
0
9 2-In XOR~
219 503 399 0 3 22
0 37 37 23
0
0 0 624 0
4 4070
-14 -24 14 -16
3 U4A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 1 2 0
1 U
3747 0 0
0
0
9 2-In XOR~
219 503 455 0 3 22
0 37 37 18
0
0 0 624 0
4 4070
-14 -24 14 -16
3 U2D
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 4 1 0
1 U
3549 0 0
0
0
9 2-In XOR~
219 504 521 0 3 22
0 37 37 17
0
0 0 624 0
4 4070
-14 -24 14 -16
3 U2C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 3 1 0
1 U
7931 0 0
0
0
9 2-In XOR~
219 507 586 0 3 22
0 37 37 16
0
0 0 624 0
4 4070
-14 -24 14 -16
3 U2B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 2 1 0
1 U
9325 0 0
0
0
9 V Source~
197 68 630 0 2 5
0 30 37
0
0 0 17264 0
3 10V
13 0 34 8
3 Vs1
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
8903 0 0
0
0
12 SPDT Switch~
164 179 296 0 3 11
0 37 30 37
0
0 0 4720 0
0
2 A1
-8 -15 6 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
3834 0 0
0
0
12 SPDT Switch~
164 180 267 0 3 11
0 37 30 37
0
0 0 4720 0
0
2 A2
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
3363 0 0
0
0
12 SPDT Switch~
164 187 242 0 3 11
0 37 30 37
0
0 0 4720 0
0
2 A3
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
7668 0 0
0
0
12 SPDT Switch~
164 187 213 0 3 11
0 37 30 37
0
0 0 4720 0
0
2 A4
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
4718 0 0
0
0
12 SPDT Switch~
164 182 183 0 3 11
0 37 30 37
0
0 0 4720 0
0
2 A5
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
3874 0 0
0
0
12 SPDT Switch~
164 185 156 0 3 11
0 37 30 37
0
0 0 4720 0
0
2 A6
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
6671 0 0
0
0
12 SPDT Switch~
164 186 125 0 3 11
0 37 30 37
0
0 0 4720 0
0
2 A7
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
3789 0 0
0
0
12 SPDT Switch~
164 184 95 0 3 11
0 37 30 37
0
0 0 4720 0
0
2 A8
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
4871 0 0
0
0
12 SPDT Switch~
164 185 558 0 3 11
0 37 30 37
0
0 0 4720 0
0
2 B2
-8 -16 6 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
3750 0 0
0
0
12 SPDT Switch~
164 184 529 0 3 11
0 37 30 37
0
0 0 4720 0
0
2 B3
-8 -16 6 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
8778 0 0
0
0
12 SPDT Switch~
164 183 503 0 3 11
0 37 30 37
0
0 0 4720 0
0
2 B4
-8 -16 6 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
538 0 0
0
0
12 SPDT Switch~
164 183 476 0 3 11
0 37 30 37
0
0 0 4720 0
0
2 B5
-8 -16 6 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
6843 0 0
0
0
12 SPDT Switch~
164 181 447 0 3 11
0 37 30 37
0
0 0 4720 0
0
2 B6
-8 -16 6 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
3136 0 0
0
0
12 SPDT Switch~
164 183 419 0 3 11
0 37 30 37
0
0 0 4720 0
0
2 B7
-8 -16 6 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
5950 0 0
0
0
12 SPDT Switch~
164 182 391 0 3 11
0 37 30 37
0
0 0 4720 0
0
2 B8
-8 -16 6 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
5670 0 0
0
0
12 SPDT Switch~
164 184 591 0 10 11
0 30 30 37 0 0 0 0 0 0
1
0
0 0 4720 0
0
2 B1
-8 -16 6 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
6828 0 0
0
0
9 2-In XOR~
219 506 639 0 3 22
0 37 30 15
0
0 0 624 0
4 4070
-14 -24 14 -16
3 U2A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 1096765229
65 0 0 0 4 1 1 0
1 U
6735 0 0
0
0
7 Ground~
168 120 670 0 1 3
0 37
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8365 0 0
0
0
9 Resistor~
219 867 626 0 3 5
0 37 28 -1
0
0 0 880 90
3 300
5 0 26 8
2 R9
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4132 0 0
0
0
9 Resistor~
219 924 631 0 3 5
0 37 3 -1
0
0 0 880 90
3 300
5 0 26 8
2 R8
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4551 0 0
0
0
9 Resistor~
219 960 632 0 3 5
0 37 4 -1
0
0 0 880 90
3 300
5 0 26 8
2 R7
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3635 0 0
0
0
9 Resistor~
219 995 634 0 3 5
0 37 5 -1
0
0 0 880 90
3 300
5 0 26 8
2 R6
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3973 0 0
0
0
9 Resistor~
219 1032 630 0 3 5
0 37 9 -1
0
0 0 880 90
3 300
5 0 26 8
2 R5
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3851 0 0
0
0
9 Resistor~
219 1070 629 0 3 5
0 37 6 -1
0
0 0 880 90
3 300
5 0 26 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8383 0 0
0
0
9 Resistor~
219 1111 631 0 3 5
0 37 7 -1
0
0 0 880 90
3 300
5 0 26 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9334 0 0
0
0
9 Resistor~
219 1151 633 0 3 5
0 37 8 -1
0
0 0 880 90
3 300
5 0 26 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7471 0 0
0
0
9 Resistor~
219 1191 634 0 3 5
0 37 10 -1
0
0 0 880 90
3 300
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3334 0 0
0
0
89
1 0 37 0 0 0 2 1 0 0 47 2
145 348
145 348
1 1 37 0 0 8320 2 31 0 0 57 3
867 644
867 664
120 664
1 0 37 0 0 0 2 32 0 0 10 2
924 649
924 664
1 0 37 0 0 0 2 33 0 0 10 2
960 650
960 664
1 0 37 0 0 0 2 34 0 0 10 2
995 652
995 664
1 0 37 0 0 0 2 35 0 0 10 2
1032 648
1032 664
1 0 37 0 0 0 2 36 0 0 10 2
1070 647
1070 664
1 0 37 0 0 0 2 37 0 0 10 2
1111 649
1111 664
1 0 37 0 0 0 2 38 0 0 10 2
1151 651
1151 664
1 0 37 0 0 0 2 39 0 0 2 3
1191 652
1191 664
867 664
10 2 3 0 0 8320 0 3 32 0 0 3
848 443
924 443
924 613
11 2 4 0 0 8320 0 3 33 0 0 3
848 452
960 452
960 614
12 2 5 0 0 8320 0 3 34 0 0 3
848 461
995 461
995 616
10 2 6 0 0 8320 0 2 36 0 0 3
840 168
1070 168
1070 611
11 2 7 0 0 8320 0 2 37 0 0 3
840 177
1111 177
1111 613
12 2 8 0 0 8320 0 2 38 0 0 3
840 186
1151 186
1151 615
13 2 9 0 0 4224 0 3 35 0 0 3
848 470
1032 470
1032 612
13 2 10 0 0 8320 0 2 39 0 0 3
840 195
1191 195
1191 616
3 0 37 0 0 0 2 25 0 0 57 2
164 451
125 451
1 1 37 0 0 4224 11 20 3 0 0 4
201 95
741 95
741 416
784 416
2 1 37 0 0 12416 12 3 19 0 0 6
784 425
725 425
725 107
221 107
221 125
203 125
3 1 37 0 0 12416 13 3 18 0 0 6
784 434
711 434
711 120
236 120
236 156
202 156
4 1 37 0 0 12416 14 3 17 0 0 6
784 443
699 443
699 131
249 131
249 183
199 183
3 8 15 0 0 8320 0 29 2 0 0 4
539 639
644 639
644 204
776 204
7 3 16 0 0 8320 0 2 11 0 0 4
776 195
631 195
631 586
540 586
3 6 17 0 0 8320 0 10 2 0 0 4
537 521
618 521
618 186
776 186
5 3 18 0 0 8320 0 2 9 0 0 6
776 177
606 177
606 439
547 439
547 455
536 455
1 1 37 0 0 4224 19 2 16 0 0 4
776 141
262 141
262 213
204 213
2 1 37 0 0 4224 20 2 15 0 0 4
776 150
286 150
286 242
204 242
3 1 37 0 0 4224 21 2 14 0 0 4
776 159
311 159
311 267
197 267
4 1 37 0 0 4224 22 2 13 0 0 4
776 168
331 168
331 296
196 296
8 3 23 0 0 4224 0 3 8 0 0 4
784 479
560 479
560 399
536 399
7 3 24 0 0 4224 0 3 7 0 0 4
784 470
572 470
572 319
536 319
6 3 25 0 0 4224 0 3 6 0 0 4
784 461
583 461
583 268
532 268
5 3 26 0 0 8320 0 3 5 0 0 4
784 452
593 452
593 214
534 214
0 9 37 0 0 4224 27 0 2 53 0 4
437 344
686 344
686 222
776 222
14 2 28 0 0 8320 0 3 31 0 0 3
848 497
867 497
867 608
14 9 29 0 0 12416 0 2 3 0 0 6
840 222
852 222
852 377
685 377
685 497
784 497
2 1 30 0 0 12416 0 29 28 0 0 4
490 648
400 648
400 591
201 591
2 1 37 0 0 12416 31 11 21 0 0 4
491 595
416 595
416 558
202 558
2 1 37 0 0 8320 32 10 22 0 0 3
488 530
488 529
201 529
2 1 37 0 0 12416 33 9 23 0 0 4
487 464
415 464
415 503
200 503
2 1 37 0 0 12416 34 8 24 0 0 4
487 408
397 408
397 476
200 476
2 1 37 0 0 12416 35 7 25 0 0 4
487 328
380 328
380 447
198 447
2 1 37 0 0 12416 36 6 26 0 0 4
483 277
364 277
364 419
200 419
1 2 37 0 0 8320 0 27 5 0 0 4
199 391
351 391
351 223
485 223
3 0 37 0 0 0 2 4 0 0 82 2
271 348
125 348
0 2 30 0 0 4096 38 0 4 71 0 3
68 339
271 339
271 340
0 1 37 0 0 0 27 0 29 50 0 3
437 577
437 630
490 630
1 0 37 0 0 0 27 11 0 0 51 3
491 577
437 577
437 512
1 0 37 0 0 0 27 10 0 0 52 3
488 512
437 512
437 446
1 0 37 0 0 0 27 9 0 0 53 3
487 446
437 446
437 390
1 0 37 0 0 0 27 8 0 0 56 3
487 390
437 390
437 344
1 0 37 0 0 0 27 7 0 0 56 2
487 310
437 310
1 0 37 0 0 0 27 6 0 0 56 2
483 259
437 259
1 1 37 0 0 0 27 5 4 0 0 4
485 205
437 205
437 344
305 344
0 1 37 0 0 128 2 0 30 0 0 3
125 375
125 664
120 664
3 0 37 0 0 0 2 28 0 0 57 2
167 595
125 595
3 0 37 0 0 0 2 21 0 0 57 2
168 562
125 562
3 0 37 0 0 0 2 22 0 0 57 2
167 533
125 533
3 0 37 0 0 0 2 23 0 0 57 2
166 507
125 507
3 0 37 0 0 0 2 24 0 0 57 2
166 480
125 480
3 0 37 0 0 0 2 26 0 0 57 2
166 423
125 423
3 0 37 0 0 0 2 27 0 0 57 2
165 395
125 395
2 0 30 0 0 0 38 27 0 0 71 2
165 387
68 387
2 0 30 0 0 0 38 26 0 0 71 2
166 415
68 415
2 0 30 0 0 0 38 25 0 0 71 2
164 443
68 443
2 0 30 0 0 0 38 24 0 0 71 2
166 472
68 472
2 0 30 0 0 0 38 23 0 0 71 2
166 499
68 499
2 0 30 0 0 0 38 22 0 0 71 2
167 525
68 525
2 2 30 0 0 8320 38 21 20 0 0 4
168 554
68 554
68 91
167 91
2 0 30 0 0 0 38 28 0 0 74 2
167 587
68 587
1 2 37 0 0 0 2 30 12 0 0 3
120 664
68 664
68 651
1 0 30 0 0 0 38 12 0 0 71 3
68 609
68 554
69 554
3 0 37 0 0 0 2 13 0 0 82 2
162 300
125 300
3 0 37 0 0 0 2 14 0 0 82 2
163 271
125 271
3 0 37 0 0 0 2 15 0 0 82 2
170 246
125 246
3 0 37 0 0 0 2 16 0 0 82 2
170 217
125 217
3 0 37 0 0 0 2 17 0 0 82 2
165 187
125 187
3 0 37 0 0 0 2 18 0 0 82 2
168 160
125 160
3 0 37 0 0 0 2 19 0 0 82 2
169 129
125 129
3 0 37 0 0 128 2 20 0 0 0 3
167 99
125 99
125 376
2 0 30 0 0 0 38 13 0 0 71 2
162 292
68 292
2 0 30 0 0 0 38 14 0 0 71 2
163 263
68 263
2 0 30 0 0 0 38 15 0 0 71 2
170 238
68 238
2 0 30 0 0 0 38 16 0 0 71 2
170 209
68 209
2 0 30 0 0 0 38 17 0 0 71 2
165 179
68 179
2 0 30 0 0 0 38 18 0 0 71 2
168 152
68 152
2 0 30 0 0 0 38 19 0 0 71 2
169 121
68 121
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
1312660 1210432 100 100 0 0
0 0 0 0
1 66 162 136
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12401 0
4 2 2
1
791 284
0 11 0 0 2	0 90 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
