CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
0 66 1280 980
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 66 1280 980
144179218 0
0
6 Title:
5 Name:
0
0
0
50
12 SPST Switch~
165 833 32 0 10 11
0 17 17 0 0 0 0 0 0 0
1
0
0 0 4720 0
0
3 S13
-11 -18 10 -10
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
8953 0 0
0
0
12 SPST Switch~
165 795 715 0 10 11
0 18 18 0 0 0 0 0 0 0
1
0
0 0 4720 0
0
3 S12
-11 -18 10 -10
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
4441 0 0
0
0
12 SPST Switch~
165 74 435 0 10 11
0 18 18 0 0 0 0 0 0 0
1
0
0 0 4720 90
0
3 S11
10 -6 31 2
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
3618 0 0
0
0
12 SPST Switch~
165 76 196 0 10 11
0 12 12 0 0 0 0 0 0 0
1
0
0 0 4720 90
0
3 S10
10 -6 31 2
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
6153 0 0
0
0
11 Multimeter~
205 846 320 0 21 21
0 17 23 24 18 0 0 0 0 0
32 50 52 46 48 48 77 101 0 0
4 73
0
0 0 16464 270
6 1.000u
-21 -37 21 -29
3 MM1
-11 -47 10 -39
0
0
31 R1%D %1 %2 1E-9
%D %4 %2 DC %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
73 0 0 0 0 0 0 0
1 I
5394 0 0
0
0
12 SPST Switch~
165 193 282 0 2 11
0 10 8
0
0 0 4720 90
0
2 S9
11 -6 25 2
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
7734 0 0
0
0
12 SPST Switch~
165 286 259 0 10 11
0 10 10 0 0 0 0 0 0 0
1
0
0 0 4720 0
0
2 S8
-7 -18 7 -10
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
9914 0 0
0
0
12 SPST Switch~
165 214 84 0 10 11
0 12 12 0 0 0 0 0 0 0
1
0
0 0 4720 90
0
2 S6
11 -6 25 2
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3747 0 0
0
0
12 SPST Switch~
165 243 67 0 2 11
0 13 12
0
0 0 4720 0
0
2 S7
-7 -41 7 -33
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3549 0 0
0
0
12 SPST Switch~
165 596 290 0 2 11
0 5 15
0
0 0 4720 90
0
2 S5
11 -6 25 2
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
7931 0 0
0
0
12 SPST Switch~
165 572 268 0 10 11
0 5 5 0 0 0 0 0 0 0
1
0
0 0 4720 0
0
2 S4
-7 -18 7 -10
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
9325 0 0
0
0
12 SPST Switch~
165 993 406 0 10 11
0 18 18 0 0 0 0 0 0 0
1
0
0 0 4720 90
0
2 S3
11 -6 25 2
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
8903 0 0
0
0
12 SPST Switch~
165 962 192 0 10 11
0 17 17 0 0 0 0 0 0 0
1
0
0 0 4720 0
0
2 S2
-7 -18 7 -10
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3834 0 0
0
0
12 SPST Switch~
165 905 211 0 2 11
0 17 19
0
0 0 4720 90
0
2 S1
11 -6 25 2
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3363 0 0
0
0
11 Multimeter~
205 267 328 0 21 21
0 10 25 26 9 0 0 0 0 0
32 55 46 48 49 56 32 86 0 0
0 82
0
0 0 16464 270
8 100.0Meg
-28 -36 28 -28
4 MM10
-14 -46 14 -38
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
1 R
7668 0 0
0
0
11 Multimeter~
205 176 227 0 21 21
0 14 27 28 10 0 0 0 0 0
32 49 57 46 48 50 109 65 0 0
0 86
0
0 0 16464 782
6 1.000u
-21 -36 21 -28
3 MM9
-11 -46 10 -38
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 1 0 0 0
1 V
4718 0 0
0
0
11 Multimeter~
205 1215 258 0 21 21
0 17 29 30 18 0 0 0 0 0
32 50 52 46 48 48 32 86 0 0
0 82
0
0 0 16464 270
8 100.0Meg
-28 -36 28 -28
3 MM8
-11 -46 10 -38
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
1 R
3874 0 0
0
0
11 Multimeter~
205 111 116 0 21 21
0 12 31 32 14 0 0 0 0 0
32 49 50 46 48 55 32 86 0 0
0 82
0
0 0 16464 782
8 100.0Meg
-28 -36 28 -28
3 MM7
-11 -46 10 -38
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
1 R
6671 0 0
0
0
11 Multimeter~
205 524 442 0 21 21
0 22 33 34 18 0 0 0 0 0
32 52 46 57 49 53 32 86 0 0
0 82
0
0 0 16464 270
8 100.0Meg
-28 -36 28 -28
3 MM6
-11 -46 10 -38
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
1 R
3789 0 0
0
0
11 Multimeter~
205 705 329 0 21 21
0 5 35 36 18 0 0 0 0 0
32 49 49 46 57 51 32 86 0 0
0 82
0
0 0 16464 270
8 100.0Meg
-28 -36 28 -28
3 MM4
-11 -46 10 -38
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
1 R
4871 0 0
0
0
11 Multimeter~
205 49 313 0 21 21
0 12 37 38 18 0 0 0 0 0
32 50 52 46 48 48 32 86 0 0
0 82
0
0 0 16464 782
8 100.0Meg
-28 -36 28 -28
3 MM3
-11 -46 10 -38
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
1 R
3750 0 0
0
0
11 Multimeter~
205 310 403 0 21 21
0 9 39 40 22 0 0 0 0 0
32 49 49 46 49 50 109 65 0 0
0 86
0
0 0 16464 0
6 1.000u
-21 -19 21 -11
3 MM2
-11 -29 10 -21
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 1 0 0 0
1 V
8778 0 0
0
0
11 Multimeter~
205 476 187 0 21 21
0 14 41 42 5 0 0 0 0 0
32 52 49 46 52 51 109 65 0 0
0 86
0
0 0 16464 0
6 1.000u
-21 -19 21 -11
3 MM1
-11 -29 10 -21
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 1 0 0 0
1 V
538 0 0
0
0
11 Multimeter~
205 678 9 0 21 21
0 12 43 44 17 0 0 0 0 0
32 50 54 46 54 54 109 65 0 0
0 86
0
0 0 16464 0
6 1.000u
-21 -19 21 -11
3 MM0
-11 -29 10 -21
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 1 0 0 0
1 V
6843 0 0
0
0
7 Ground~
168 127 764 0 1 3
0 18
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3136 0 0
0
0
9 V Source~
197 76 318 0 2 5
0 12 18
0
0 0 17264 0
3 24V
13 0 34 8
3 Vs1
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
5950 0 0
0
0
9 Resistor~
219 432 309 0 2 5
0 9 10
0
0 0 880 90
3 369
8 0 29 8
3 R24
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
5670 0 0
0
0
9 Resistor~
219 437 137 0 2 5
0 14 13
0
0 0 880 90
3 198
8 0 29 8
3 R23
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
6828 0 0
0
0
9 Resistor~
219 513 322 0 3 5
0 18 5 -1
0
0 0 880 90
3 288
8 0 29 8
3 R22
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
6735 0 0
0
0
9 Resistor~
219 891 337 0 2 5
0 18 19
0
0 0 880 90
3 900
8 1 29 9
3 R21
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
8365 0 0
0
0
9 Resistor~
219 337 127 0 2 5
0 14 12
0
0 0 880 90
5 1.25k
1 0 36 8
3 R20
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4132 0 0
0
0
9 Resistor~
219 302 127 0 2 5
0 14 12
0
0 0 880 90
5 1.15k
1 0 36 8
3 R19
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4551 0 0
0
0
9 Resistor~
219 268 126 0 2 5
0 14 12
0
0 0 880 90
5 1.15k
1 0 36 8
3 R18
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3635 0 0
0
0
9 Resistor~
219 235 125 0 2 5
0 14 12
0
0 0 880 90
5 1.15k
1 0 36 8
3 R17
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3973 0 0
0
0
9 Resistor~
219 204 125 0 2 5
0 14 12
0
0 0 880 90
5 1.07k
1 0 36 8
3 R16
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3851 0 0
0
0
9 Resistor~
219 172 123 0 2 5
0 14 12
0
0 0 880 90
4 1.5k
4 0 32 8
3 R11
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8383 0 0
0
0
9 Resistor~
219 149 326 0 2 5
0 9 8
0
0 0 880 90
3 750
7 0 28 8
3 R15
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
9334 0 0
0
0
9 Resistor~
219 644 334 0 3 5
0 18 15 -1
0
0 0 880 90
5 1.18k
2 0 37 8
3 R10
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
7471 0 0
0
0
9 Resistor~
219 615 335 0 3 5
0 18 15 -1
0
0 0 880 90
5 1.15k
-2 0 33 8
2 R9
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
3334 0 0
0
0
9 Resistor~
219 587 333 0 3 5
0 18 15 -1
0
0 0 880 90
5 1.15k
-2 0 33 8
2 R8
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
3559 0 0
0
0
9 Resistor~
219 558 333 0 3 5
0 18 15 -1
0
0 0 880 90
5 1.15k
-2 0 33 8
2 R7
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
984 0 0
0
0
9 Resistor~
219 1110 340 0 2 5
0 18 17
0
0 0 880 90
5 5.49k
-2 0 33 8
2 R6
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
7557 0 0
0
0
9 Resistor~
219 1078 340 0 2 5
0 18 17
0
0 0 880 90
5 5.49k
-2 0 33 8
2 R5
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
3146 0 0
0
0
9 Resistor~
219 1044 337 0 2 5
0 18 17
0
0 0 880 90
5 5.36k
-2 0 33 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
5687 0 0
0
0
9 Resistor~
219 1009 336 0 2 5
0 18 17
0
0 0 880 90
5 5.36k
-2 0 33 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
7939 0 0
0
0
9 Resistor~
219 975 336 0 2 5
0 18 17
0
0 0 880 90
5 5.36k
-2 0 33 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
3308 0 0
0
0
9 Resistor~
219 942 336 0 2 5
0 18 17
0
0 0 880 90
5 5.36k
-2 0 33 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
3408 0 0
0
0
9 Resistor~
219 412 443 0 3 5
0 18 22 -1
0
0 0 880 90
3 442
8 0 29 8
3 R14
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9773 0 0
0
0
9 Resistor~
219 195 535 0 3 5
0 18 9 -1
0
0 0 880 90
3 622
8 0 29 8
3 R13
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
691 0 0
0
0
9 Resistor~
219 193 324 0 2 5
0 9 8
0
0 0 880 90
3 732
8 0 29 8
3 R12
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7834 0 0
0
0
88
1 0 17 0 0 4224 3 1 0 0 8 2
850 32
891 32
1 0 18 0 0 12416 4 2 0 0 31 4
812 715
812 714
917 714
917 527
4 0 18 0 0 0 4 5 0 0 27 3
830 352
830 498
917 498
1 0 17 0 0 4096 3 5 0 0 8 3
830 302
830 153
906 153
0 0 18 0 0 4224 2 0 0 58 74 3
600 353
600 714
412 714
0 1 5 0 0 4224 0 0 10 0 0 2
597 249
597 272
0 2 18 0 0 128 2 0 2 5 0 3
600 714
778 714
778 715
0 1 17 0 0 12288 3 0 14 0 0 4
887 33
887 32
906 32
906 193
2 0 18 0 0 0 2 3 0 0 82 3
75 451
75 715
127 715
2 1 12 0 0 8336 6 4 26 0 0 3
77 212
76 212
76 297
1 0 10 0 0 8192 7 15 0 0 15 3
251 310
232 310
232 259
2 2 8 0 0 8192 0 6 50 0 0 3
194 298
193 298
193 306
1 0 9 0 0 8320 0 27 0 0 87 3
432 327
432 382
195 382
1 2 10 0 0 4224 0 7 27 0 0 3
303 259
432 259
432 291
0 2 10 0 0 4224 7 0 7 53 0 2
193 259
269 259
0 2 12 0 0 8192 11 0 8 41 0 3
217 107
215 107
215 100
1 0 12 0 0 4096 0 8 0 0 21 2
215 66
215 65
0 0 12 0 0 4096 0 0 0 21 88 2
200 65
200 43
1 2 13 0 0 8320 0 9 28 0 0 4
260 67
260 68
437 68
437 119
1 0 14 0 0 8192 0 28 0 0 85 4
437 155
437 194
397 194
397 209
1 2 12 0 0 8192 0 18 9 0 0 4
127 98
127 65
226 65
226 67
2 0 15 0 0 4096 0 10 0 0 61 2
597 306
597 317
1 0 5 0 0 0 0 11 0 0 54 2
589 268
597 268
1 0 18 0 0 0 2 29 0 0 5 3
513 340
513 398
600 398
2 2 5 0 0 8320 16 29 11 0 0 3
513 304
513 268
555 268
0 1 18 0 0 0 4 0 30 27 0 4
917 455
917 411
891 411
891 355
0 0 18 0 0 0 4 0 0 2 29 2
917 527
917 455
1 0 17 0 0 8320 0 13 0 0 72 3
979 192
1009 192
1009 318
2 0 18 0 0 0 4 12 0 0 0 4
994 422
979 422
979 455
914 455
1 0 18 0 0 4096 0 12 0 0 64 4
994 388
994 367
980 367
980 354
4 0 18 0 0 8320 4 17 0 0 0 3
1199 290
1199 527
914 527
1 0 17 0 0 8320 3 17 0 0 8 3
1199 240
1199 110
906 110
1 2 17 0 0 0 3 14 13 0 0 3
906 193
906 192
945 192
2 2 19 0 0 4224 0 14 30 0 0 3
906 227
906 319
891 319
4 2 17 0 0 4224 20 24 1 0 0 2
703 32
816 32
0 0 18 0 0 0 2 0 0 37 86 2
195 642
195 573
0 0 18 0 0 0 2 0 0 0 0 3
194 639
195 639
195 709
0 0 14 0 0 4096 0 0 0 39 48 2
224 190
224 143
4 0 14 0 0 12288 0 18 0 0 85 5
127 148
144 148
144 190
236 190
236 209
2 2 12 0 0 8192 11 35 36 0 0 3
204 107
204 105
172 105
2 2 12 0 0 0 11 34 35 0 0 2
235 107
204 107
2 2 12 0 0 8192 11 33 34 0 0 3
268 108
268 107
235 107
2 2 12 0 0 8192 11 32 33 0 0 3
302 109
302 108
268 108
2 2 12 0 0 4224 11 31 32 0 0 2
337 109
302 109
1 1 14 0 0 0 0 32 31 0 0 2
302 145
337 145
1 1 14 0 0 0 0 33 32 0 0 3
268 144
268 145
302 145
1 1 14 0 0 0 0 34 33 0 0 3
235 143
235 144
268 144
1 1 14 0 0 0 0 35 34 0 0 2
204 143
235 143
1 1 14 0 0 0 0 36 35 0 0 4
172 141
193 141
193 143
204 143
2 2 8 0 0 8320 0 50 37 0 0 3
193 306
193 308
149 308
1 1 9 0 0 0 0 37 50 0 0 3
149 344
149 342
193 342
4 0 9 0 0 0 0 15 0 0 87 2
251 360
195 360
4 1 10 0 0 0 7 16 6 0 0 4
192 259
193 259
193 264
194 264
1 0 5 0 0 8192 0 20 0 0 6 3
689 311
689 268
597 268
4 0 18 0 0 0 2 20 0 0 5 3
689 361
689 398
600 398
4 0 5 0 0 4224 0 23 0 0 6 3
501 210
597 210
597 252
1 1 18 0 0 0 2 39 38 0 0 3
615 353
615 352
644 352
1 1 18 0 0 0 2 40 39 0 0 3
587 351
587 353
615 353
1 1 18 0 0 0 2 41 40 0 0 2
558 351
587 351
2 2 15 0 0 8320 0 39 38 0 0 3
615 317
615 316
644 316
2 2 15 0 0 0 0 40 39 0 0 3
587 315
587 317
615 317
2 2 15 0 0 0 0 41 40 0 0 2
558 315
587 315
1 1 18 0 0 4096 0 46 47 0 0 2
975 354
942 354
0 1 18 0 0 8320 0 0 46 65 0 3
1012 355
1012 354
975 354
1 1 18 0 0 0 0 45 44 0 0 3
1009 354
1009 355
1044 355
0 1 18 0 0 0 0 0 44 67 0 3
1060 358
1044 358
1044 355
1 0 18 0 0 0 0 43 0 0 0 2
1078 358
1060 358
1 1 18 0 0 0 0 42 43 0 0 2
1110 358
1078 358
2 2 17 0 0 0 0 43 42 0 0 2
1078 322
1110 322
2 2 17 0 0 0 0 44 43 0 0 3
1044 319
1044 322
1078 322
2 2 17 0 0 0 0 45 44 0 0 3
1009 318
1009 319
1044 319
2 2 17 0 0 0 0 46 45 0 0 2
975 318
1009 318
2 2 17 0 0 0 0 47 46 0 0 2
942 318
975 318
0 0 18 0 0 0 2 0 0 83 75 3
412 705
412 715
195 715
0 0 18 0 0 0 2 0 0 37 9 3
195 703
195 715
127 715
0 1 18 0 0 4096 21 0 3 78 0 2
75 380
75 417
1 0 12 0 0 0 6 21 0 0 10 3
65 295
65 229
76 229
4 2 18 0 0 12416 21 21 26 0 0 4
65 345
65 380
76 380
76 339
4 0 18 0 0 0 2 19 0 0 83 4
508 474
427 474
427 475
412 475
1 2 22 0 0 4224 0 19 48 0 0 4
508 424
427 424
427 425
412 425
4 2 22 0 0 0 0 22 48 0 0 3
335 426
335 425
412 425
1 0 18 0 0 0 2 25 0 0 0 2
127 758
127 709
1 0 18 0 0 0 2 48 0 0 0 2
412 461
412 709
0 1 9 0 0 0 0 0 22 87 0 3
195 425
285 425
285 426
1 1 14 0 0 4224 0 16 23 0 0 3
192 209
451 209
451 210
1 0 18 0 0 0 2 49 0 0 0 3
195 553
195 589
194 589
1 2 9 0 0 0 0 50 49 0 0 3
193 342
195 342
195 517
1 1 12 0 0 8336 0 24 4 0 0 5
653 32
653 43
76 43
76 178
77 178
10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
905 277 985 301
915 285 987 301
9 Req = 900
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
504 278 584 302
514 286 586 302
9 Req = 288
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
708 26 772 50
718 34 774 50
7 26.7 mA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
509 182 573 206
519 190 575 206
7 41.7 mA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
338 399 402 423
348 407 404 423
7 12.0 mA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
415 483 551 507
425 491 553 507
16 V=4.95 to 5.05 V
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
715 308 827 352
725 316 829 348
22 V = 11.88 to 
12.12V
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
1075 223 1163 267
1085 231 1165 263
22 V = 23.76 
to 24.24V
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
346 262 426 286
356 269 428 285
9 Req = 369
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
448 92 528 116
458 100 530 116
9 Req = 197
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 1e-006 1e-007 1e-007
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
3278160 1079360 100 100 0 0
0 0 0 0
558 222 719 292
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12401 0
4 5 10
1
306 209
0 14 0 0 1	0 85 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
