CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 120 9
32 88 1248 734
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
32 88 1248 734
144179218 256
0
6 Title:
5 Name:
0
0
0
4
7 Ground~
168 162 324 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8953 0 0
0
0
6 Diode~
219 378 270 0 2 5
0 4 2
0
0 0 1616 270
5 DIODE
17 0 52 8
4 Vout
15 -10 43 -2
18 Channel B / Output
-127 29 -1 37
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
4441 0 0
0
0
4 VCO~
221 189 243 0 5 9
0 3 2 3 2 3
0
0 0 1616 0
6 TRIVCO
37 -2 79 6
3 Vs1
-18 -28 3 -20
18 Channel A and Sync
32 -18 158 -10
0
29 %D %%vd(%1,%2) %%vd(%3,%4) %M
0
13 alias:ATRIVCO
0
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 0 0 0 0
1 V
3618 0 0
0
0
9 Resistor~
219 306 189 0 2 5
0 3 4
0
0 0 880 0
3 10k
-10 -14 11 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6153 0 0
0
0
6
1 0 0 0 0 0 0 1 0 0 4 4
162 318
162 327
162 327
162 318
4 0 2 0 0 4096 0 3 0 0 4 2
198 273
198 318
3 0 3 0 0 4096 0 3 0 0 6 2
198 219
198 189
2 2 2 0 0 8320 0 2 3 0 0 4
378 280
378 318
162 318
162 273
2 1 4 0 0 8320 0 4 2 0 0 3
324 189
378 189
378 260
1 1 3 0 0 8320 0 3 4 0 0 3
162 219
162 189
288 189
2
13 7 0 0 0 0 0 0 0 0 0 0 54
11 Ubuntu Mono
0 0 0 1
359 275 373 292
362 277 369 290
1 -
13 7 0 0 0 0 0 0 0 0 0 0 54
11 Ubuntu Mono
0 0 0 1
361 234 375 251
364 236 371 249
1 +
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
524572 1210432 100 100 0 0
0 0 0 0
1 58 139 113
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12401 0
4 0.3 0.5
1
198 203
0 3 0 0 1	0 3 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
