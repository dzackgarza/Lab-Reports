CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
30 50 30 200 9
0 67 1280 765
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 67 1280 765
211288082 256
0
6 Title:
5 Name:
0
0
0
8
11 Multimeter~
205 324 81 0 21 21
0 6 7 8 5 0 0 0 0 0
45 51 57 46 49 50 110 65 0 0
0 86
0
0 0 16464 512
6 1.000u
-21 -19 21 -11
3 MM1
-11 -29 10 -21
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 0 0 0 0
1 V
8953 0 0
0
0
11 Multimeter~
205 243 126 0 21 21
0 5 9 10 3 0 0 0 0 0
45 50 48 48 46 48 117 65 0 0
0 86
0
0 0 16464 782
6 1.000u
-21 -19 21 -11
3 MM3
-11 -29 10 -21
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 1 0 0 0
1 V
4441 0 0
0
0
11 Multimeter~
205 414 81 0 21 21
0 4 11 12 6 0 0 0 0 0
45 52 46 48 48 48 32 86 0 0
0 82
0
0 0 16464 512
8 100.0Meg
-28 -19 28 -11
3 MM1
-11 -29 10 -21
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
1 R
3618 0 0
0
0
11 Multimeter~
205 207 216 0 21 21
0 3 13 14 2 0 0 0 0 0
32 49 48 46 48 48 32 86 0 0
0 82
0
0 0 16464 782
8 100.0Meg
-28 -36 28 -28
3 MM0
-11 -46 10 -38
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
1 R
6153 0 0
0
0
7 Ground~
168 264 313 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5394 0 0
0
0
9 V Source~
197 264 220 0 2 5
0 3 2
0
0 0 17136 0
2 10
16 0 30 8
3 Vs1
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
7734 0 0
0
0
9 Resistor~
219 534 221 0 3 5
0 2 4 -1
0
0 0 880 90
3 30k
19 2 40 10
2 R2
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9914 0 0
0
0
9 Resistor~
219 382 162 0 2 5
0 5 4
0
0 0 880 692
3 20k
-11 -14 10 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3747 0 0
0
0
10
1 1 3 0 0 8320 0 4 6 0 0 3
223 198
223 199
264 199
4 0 2 0 0 4096 0 4 0 0 8 2
223 248
264 248
2 0 4 0 0 4224 0 8 0 0 4 3
400 162
479 162
479 136
1 2 4 0 0 0 0 3 7 0 0 6
439 104
479 104
479 136
535 136
535 203
534 203
0 1 5 0 0 8320 0 0 8 7 0 3
299 126
299 162
364 162
1 4 6 0 0 4224 0 1 3 0 0 2
349 104
389 104
1 4 5 0 0 0 0 2 1 0 0 5
259 108
270 108
270 126
299 126
299 104
2 0 2 0 0 4096 0 6 0 0 10 2
264 241
264 283
4 1 3 0 0 128 0 2 6 0 0 3
259 158
264 158
264 199
1 1 2 0 0 8336 0 5 7 0 0 4
264 307
264 282
534 282
534 239
4
13 7 0 0 0 0 0 0 0 0 0 0 54
11 Ubuntu Mono
0 0 0 12
269 55 360 72
272 57 356 70
12 I(Voltmeter)
13 7 0 0 0 0 0 0 0 0 0 0 54
11 Ubuntu Mono
0 0 0 9
383 55 453 72
386 57 449 70
9 Voltmeter
13 7 0 0 0 0 0 0 0 0 0 0 54
11 Ubuntu Mono
0 0 0 5
166 117 208 134
169 119 204 132
5 I(s1)
13 7 0 0 0 0 0 0 0 0 0 0 54
11 Ubuntu Mono
0 0 0 15
419 180 531 197
422 182 527 195
15 Varied Resistor
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 1e-006 1e-007 1e-007
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
3736020 1210432 100 100 0 0
0 0 0 0
1 58 139 113
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 3 5
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
