CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
30 50 30 200 9
0 67 1305 765
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 67 1305 765
211288082 256
0
6 Title:
5 Name:
0
0
0
8
11 Multimeter~
205 477 180 0 21 21
0 3 7 8 4 0 0 0 0 0
78 79 32 68 65 84 65 32 0 0
0 86
0
0 0 16464 90
6 1.000u
-21 -37 21 -29
3 MM1
-11 -47 10 -39
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 0 0 0 0
1 V
8953 0 0
0
0
11 Multimeter~
205 333 117 0 21 21
0 6 9 10 5 0 0 0 0 0
78 79 32 68 65 84 65 32 0 0
0 86
0
0 0 16464 0
6 1.000u
-21 -19 21 -11
3 MM0
-11 -29 10 -21
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 0 0 0 0
1 V
4441 0 0
0
0
11 Multimeter~
205 587 201 0 21 21
0 2 11 12 4 0 0 0 0 0
78 79 32 68 65 84 65 32 0 0
0 82
0
0 0 16464 602
8 100.0Meg
-28 -19 28 -11
3 MM1
-11 -29 10 -21
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
1 R
3618 0 0
0
0
11 Multimeter~
205 207 216 0 21 21
0 6 13 14 2 0 0 0 0 0
78 79 32 68 65 84 65 32 0 0
0 82
0
0 0 16464 782
8 100.0Meg
-28 -36 28 -28
3 MM0
-11 -46 10 -38
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
1 R
6153 0 0
0
0
7 Ground~
168 264 313 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5394 0 0
0
0
9 V Source~
197 264 220 0 2 5
0 6 2
0
0 0 17136 0
1 5
19 0 26 8
3 Vs1
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
7734 0 0
0
0
9 Resistor~
219 423 144 0 2 5
0 5 4
0
0 0 880 0
5 20.2k
-17 -14 18 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9914 0 0
0
0
9 Resistor~
219 507 239 0 3 5
0 2 3 -1
0
0 0 752 90
5 30.3k
13 2 48 10
2 R2
10 -4 24 4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3747 0 0
0
0
10
1 2 3 0 0 4224 0 1 8 0 0 3
494 211
507 211
507 221
0 4 4 0 0 4096 0 0 1 4 0 3
508 145
508 161
494 161
1 0 2 0 0 8192 0 3 0 0 10 3
570 232
570 282
506 282
4 2 4 0 0 8320 0 3 7 0 0 4
570 182
570 145
441 145
441 144
1 4 5 0 0 4224 0 7 2 0 0 3
405 144
358 144
358 140
1 1 6 0 0 4224 0 6 2 0 0 4
264 199
264 144
308 144
308 140
1 1 6 0 0 128 0 4 6 0 0 3
223 198
223 199
264 199
4 0 2 0 0 0 0 4 0 0 9 2
223 248
264 248
2 0 2 0 0 0 0 6 0 0 10 2
264 241
264 283
1 1 2 0 0 8320 0 5 8 0 0 4
264 307
264 282
507 282
507 257
5
13 7 0 0 0 0 0 0 0 0 0 0 54
11 Ubuntu Mono
0 0 0 3
183 166 226 183
189 170 225 183
3 DVM
13 7 0 0 0 0 0 0 0 0 0 0 54
11 Ubuntu Mono
0 0 0 3
571 152 614 169
577 156 613 169
3 DVM
13 7 0 0 0 0 0 0 0 0 0 0 54
11 Ubuntu Mono
0 0 0 5
415 179 458 196
421 183 457 196
5 I(R2)
13 7 0 0 0 0 0 0 0 0 0 0 54
11 Ubuntu Mono
0 0 0 15
384 230 502 247
390 234 501 247
15 Varied Resistor
13 7 0 0 0 0 0 0 0 0 0 0 54
11 Ubuntu Mono
0 0 0 5
254 110 296 127
257 112 292 125
5 I(s1)
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 1e-006 1e-007 1e-007
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
1575304 1079360 100 100 0 0
0 0 0 0
1 58 162 128
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 2e-007 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
