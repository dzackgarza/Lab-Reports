CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
210 80 30 200 9
32 89 1248 744
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
32 89 1248 744
211288082 256
0
6 Title:
5 Name:
0
0
0
7
11 Multimeter~
205 639 162 0 21 21
0 6 9 10 4 0 0 0 0 0
78 79 32 68 65 84 65 32 0 0
0 86
0
0 0 16448 270
6 1.000u
-21 -36 21 -28
3 MM2
-11 -46 10 -38
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 1 0 0 0
1 V
8953 0 0
0
0
11 Multimeter~
205 495 162 0 21 21
0 6 11 12 5 0 0 0 0 0
78 79 32 68 65 84 65 32 0 0
0 86
0
0 0 16448 270
6 1.000u
-21 -36 21 -28
3 MM1
-11 -46 10 -38
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 1 0 0 0
1 V
4441 0 0
0
0
11 Multimeter~
205 405 99 0 21 21
0 3 13 14 6 0 0 0 0 0
78 79 32 68 65 84 65 32 0 0
0 86
0
0 0 16448 0
6 1.000u
-21 -19 21 -11
3 MM0
-11 -29 10 -21
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 1 0 0 0
1 V
3618 0 0
0
0
7 Ground~
168 333 306 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6153 0 0
0
0
9 I Source~
198 333 198 0 2 5
0 2 3
0
0 0 17248 692
5 100mA
13 0 48 8
3 Is1
20 -10 41 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
73 0 0 0 1 0 0 0
2 Is
5394 0 0
0
0
9 Resistor~
219 621 234 0 3 5
0 2 4 -1
0
0 0 864 90
3 30k
5 0 26 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7734 0 0
0
0
9 Resistor~
219 477 234 0 3 5
0 2 5 -1
0
0 0 864 90
3 20k
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9914 0 0
0
0
8
4 2 4 0 0 8320 0 1 6 0 0 3
623 194
621 194
621 216
4 2 5 0 0 8320 0 2 7 0 0 3
479 194
477 194
477 216
4 1 6 0 0 8320 0 3 1 0 0 5
430 122
430 125
621 125
621 144
623 144
0 1 6 0 0 0 0 0 2 3 0 3
477 125
477 144
479 144
1 0 2 0 0 0 0 7 0 0 7 2
477 252
477 275
1 0 2 0 0 0 0 4 0 0 7 2
333 300
333 275
1 1 2 0 0 8320 0 6 5 0 0 4
621 252
621 275
333 275
333 219
2 1 3 0 0 4224 0 5 3 0 0 4
333 177
333 125
380 125
380 122
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
786774 1210432 100 100 0 0
0 0 0 0
1 58 139 113
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12401 0
4 500 1000
1
477 268
0 2 0 0 1	0 5 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
