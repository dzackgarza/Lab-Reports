CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 90 30 200 9
32 88 1248 733
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
32 88 1248 733
144179218 256
0
6 Title:
5 Name:
0
0
0
4
7 Ground~
168 252 288 0 1 3
0 0
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8953 0 0
0
0
10 Capacitor~
219 369 234 0 1 5
0 0
0
0 0 832 90
6 0.01uF
9 0 51 8
2 C2
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
4441 0 0
0
0
9 Resistor~
219 306 189 0 1 5
0 0
0
0 0 864 0
3 10k
-10 -14 11 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3618 0 0
0
0
11 Signal Gen~
195 216 234 0 19 64
0 0 0 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1176256512 0 1065353216
20
1 10000 0 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 576 0
5 -1/1V
-18 -30 17 -22
3 Vin
-10 -40 11 -32
0
0
37 %D %1 %2 DC 0 SIN(0 1 10k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
6153 0 0
0
0
4
1 0 0 0 0 0 0 1 0 0 2 2
252 282
252 281
1 2 0 0 0 0 0 2 4 0 0 4
369 243
369 281
247 281
247 239
2 2 0 0 0 0 0 3 2 0 0 3
324 189
369 189
369 225
1 1 0 0 0 0 0 4 3 0 0 3
247 229
247 189
288 189
3
13 7 0 0 0 0 0 0 0 0 0 0 54
11 Ubuntu Mono
0 0 0 4
429 226 464 243
432 228 460 241
4 Vout
13 7 0 0 0 0 0 0 0 0 0 0 54
11 Ubuntu Mono
0 0 0 1
390 271 404 288
393 273 400 286
1 -
13 7 0 0 0 0 0 0 0 0 0 0 54
11 Ubuntu Mono
0 0 0 1
386 184 400 201
389 186 396 199
1 +
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
