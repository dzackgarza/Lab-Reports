CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
20 110 30 200 9
32 88 1248 733
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
32 88 1248 733
144179218 256
0
6 Title:
5 Name:
0
0
0
6
9 Resistor~
219 414 225 0 1 5
0 0
0
0 0 864 90
2 1k
8 0 22 8
3 R5b
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8953 0 0
0
0
10 Capacitor~
219 342 180 0 1 5
0 0
0
0 0 832 180
3 1uF
-11 -18 10 -10
3 C5b
-10 -28 11 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
4441 0 0
0
0
10 Capacitor~
219 279 225 0 1 5
0 0
0
0 0 832 90
5 2.5uF
13 1 48 9
3 C5a
18 -10 39 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3618 0 0
0
0
9 Resistor~
219 216 180 0 1 5
0 0
0
0 0 864 0
3 200
-10 -14 11 -6
3 R5a
-9 -24 12 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6153 0 0
0
0
11 Signal Gen~
195 135 225 0 19 64
0 0 0 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1176256512 0 1065353216
20
1 10000 0 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 576 0
5 -1/1V
-18 -30 17 -22
3 Vin
-10 -40 11 -32
0
0
37 %D %1 %2 DC 0 SIN(0 1 10k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
5394 0 0
0
0
7 Ground~
168 189 288 0 1 3
0 0
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7734 0 0
0
0
7
1 0 0 0 0 0 0 6 0 0 3 4
189 282
189 290
189 290
189 280
1 0 0 0 0 0 0 3 0 0 3 2
279 234
279 280
1 2 0 0 0 0 0 1 5 0 0 4
414 243
414 280
166 280
166 230
2 0 0 0 0 0 0 3 0 0 6 2
279 216
279 180
1 2 0 0 0 0 0 2 1 0 0 3
351 180
414 180
414 207
2 2 0 0 0 0 0 2 4 0 0 2
333 180
234 180
1 1 0 0 0 0 0 5 4 0 0 3
166 220
166 180
198 180
3
13 7 0 0 0 0 0 0 0 0 0 0 54
11 Ubuntu Mono
0 0 0 4
449 212 484 229
452 214 480 227
4 Vout
13 7 0 0 0 0 0 0 0 0 0 0 54
11 Ubuntu Mono
0 0 0 1
428 268 442 285
431 270 438 283
1 -
13 7 0 0 0 0 0 0 0 0 0 0 54
11 Ubuntu Mono
0 0 0 1
427 178 441 195
430 180 437 193
1 +
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
