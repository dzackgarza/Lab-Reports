CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
220 90 30 400 9
32 88 1248 734
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
32 88 1248 734
144179218 256
0
6 Title:
5 Name:
0
0
0
4
10 Capacitor~
219 459 189 0 2 5
0 4 2
0
0 0 576 90
3 1uF
11 0 32 8
2 Cn
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 512 1 0 0 0
1 C
8953 0 0
0
0
9 V Source~
197 243 189 0 2 5
0 2 3
0
0 0 16992 0
3 10V
13 0 34 8
2 Vs
16 -10 30 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
4441 0 0
0
0
10 Capacitor~
219 369 189 0 2 5
0 3 2
0
0 0 576 90
3 1uF
11 0 32 8
2 C2
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3618 0 0
0
0
10 Capacitor~
219 315 189 0 2 5
0 3 2
0
0 0 576 90
3 1uF
11 0 32 8
2 C1
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6153 0 0
0
0
6
1 0 0 0 0 0 0 1 0 0 3 3
459 198
459 233
368 233
2 0 2 0 0 8320 0 1 0 0 5 3
459 180
459 126
369 126
0 1 3 0 0 4096 0 0 3 4 0 3
315 233
369 233
369 198
2 1 3 0 0 8320 0 2 4 0 0 4
243 210
243 233
315 233
315 198
0 2 2 0 0 16 0 0 3 6 0 3
315 126
369 126
369 180
1 2 2 0 0 0 0 2 4 0 0 4
243 168
243 126
315 126
315 180
1
13 7 0 0 0 0 0 0 0 0 0 0 54
11 Ubuntu Mono
0 0 0 3
411 175 439 192
414 177 435 190
3 ...
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
