CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 80 30 200 9
32 88 1248 734
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
32 88 1248 734
144179218 256
0
6 Title:
5 Name:
0
0
0
4
7 Ground~
168 216 333 0 1 3
0 0
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8953 0 0
0
0
11 Signal Gen~
195 180 252 0 19 64
0 0 0 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1176256512 0 1065353216
20
1 10000 0 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 576 0
5 -1/1V
-18 -30 17 -22
3 Vin
-10 -40 11 -32
0
0
37 %D %1 %2 DC 0 SIN(0 1 10k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
4441 0 0
0
0
9 Resistor~
219 324 252 0 1 5
0 0
0
0 0 864 90
2 1k
7 3 21 11
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3618 0 0
0
0
10 Capacitor~
219 261 207 0 1 5
0 0
0
0 0 832 0
5 100pF
-13 -18 22 -10
2 C1
-4 -28 10 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6153 0 0
0
0
4
1 0 0 0 0 0 0 1 0 0 2 4
216 327
216 332
216 332
216 320
1 2 0 0 0 0 0 3 2 0 0 4
324 270
324 320
211 320
211 257
2 2 0 0 0 0 0 4 3 0 0 3
270 207
324 207
324 234
1 1 0 0 0 0 0 2 4 0 0 3
211 247
211 207
252 207
3
13 7 0 0 0 0 0 0 0 0 0 0 54
11 Ubuntu Mono
0 0 0 4
374 246 408 262
379 248 406 260
4 Vout
13 7 0 0 0 0 0 0 0 0 0 0 54
11 Ubuntu Mono
0 0 0 1
352 302 366 318
357 304 364 316
1 -
13 7 0 0 0 0 0 0 0 0 0 0 54
11 Ubuntu Mono
0 0 0 1
348 203 362 219
353 206 360 218
1 +
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
