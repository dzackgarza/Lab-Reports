CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
20 100 30 200 9
32 88 1248 734
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
32 88 1248 734
144179218 256
0
6 Title:
5 Name:
0
0
0
6
7 Ground~
168 225 342 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8953 0 0
0
0
11 Multimeter~
205 333 234 0 17 21
0 4 6 7 3 0 0 0 0 0
78 79 32 68 65 84 65 32
0
0 0 16464 270
8 100.0Meg
-28 -36 28 -28
3 MM1
-11 -46 10 -38
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
1 R
4441 0 0
0
0
11 Multimeter~
205 270 333 0 17 21
0 3 8 9 2 0 0 0 0 0
78 79 32 68 65 84 65 32
0
0 0 16464 180
6 1.000u
-22 -19 20 -11
3 MM0
-12 -29 9 -21
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 0 0 0 0
1 V
3618 0 0
0
0
9 V Source~
197 225 261 0 2 5
0 5 2
0
0 0 17264 0
3 17V
13 0 34 8
2 Vs
16 -10 30 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
6153 0 0
0
0
9 Resistor~
219 378 243 0 2 5
0 3 4
0
0 0 624 90
2 1k
8 0 22 8
2 RL
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5394 0 0
0
0
9 Resistor~
219 225 207 0 2 5
0 5 4
0
0 0 624 90
2 1k
8 0 22 8
1 r
11 -10 18 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7734 0 0
0
0
7
0 1 2 0 0 4096 0 0 1 4 0 2
225 324
225 336
4 0 3 0 0 4096 0 2 0 0 3 2
317 266
317 324
1 1 3 0 0 4224 0 3 5 0 0 3
293 324
378 324
378 261
2 4 2 0 0 4224 0 4 3 0 0 3
225 282
225 324
243 324
1 0 4 0 0 4112 0 2 0 0 6 2
317 216
317 160
2 2 4 0 0 8320 0 6 5 0 0 4
225 189
225 160
378 160
378 225
1 1 5 0 0 4224 0 4 6 0 0 2
225 240
225 225
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
