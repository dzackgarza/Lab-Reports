CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
-3 76 997 725
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
-3 76 997 725
144179218 272
0
6 Title:
5 Name:
0
0
0
8
9 V Source~
197 57 166 0 2 5
0 5 2
0
0 0 17264 0
3 24V
13 0 34 8
2 Vs
16 -10 30 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
8953 0 0
0
0
7 Ground~
168 57 472 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4441 0 0
0
0
9 Resistor~
219 255 103 0 2 5
0 3 5
0
0 0 880 90
3 197
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3618 0 0
0
0
9 Resistor~
219 255 202 0 2 5
0 4 3
0
0 0 880 90
3 369
5 0 26 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6153 0 0
0
0
9 Resistor~
219 255 310 0 3 5
0 2 4 -1
0
0 0 880 90
3 622
5 0 26 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5394 0 0
0
0
9 Resistor~
219 624 121 0 3 5
0 2 5 -1
0
0 0 880 90
3 900
9 0 30 8
5 Load1
10 -14 45 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7734 0 0
0
0
9 Resistor~
219 489 310 0 3 5
0 2 3 -1
0
0 0 880 90
3 288
8 0 29 8
5 Load2
8 -11 43 -3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9914 0 0
0
0
9 Resistor~
219 381 310 0 3 5
0 2 4 -1
0
0 0 880 90
3 442
5 0 26 8
5 Load3
7 -10 42 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3747 0 0
0
0
11
2 0 3 0 0 8320 0 7 0 0 9 3
489 292
489 157
255 157
2 0 4 0 0 8320 0 8 0 0 8 3
381 292
381 262
255 262
1 0 2 0 0 4096 0 5 0 0 6 2
255 328
255 446
1 0 2 0 0 0 0 7 0 0 6 2
489 328
489 446
1 0 2 0 0 0 0 8 0 0 6 4
381 328
381 339
382 339
382 446
1 1 2 0 0 8320 0 2 6 0 0 4
57 466
57 446
624 446
624 139
2 1 2 0 0 0 0 1 2 0 0 2
57 187
57 466
2 1 4 0 0 0 0 5 4 0 0 2
255 292
255 220
2 1 3 0 0 0 0 4 3 0 0 2
255 184
255 121
2 0 5 0 0 4096 0 3 0 0 11 2
255 85
255 38
2 1 5 0 0 8320 0 6 1 0 0 5
624 103
624 38
56 38
56 145
57 145
12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
163 84 235 108
173 92 237 108
8 60.85 mA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
168 180 240 204
178 188 242 204
8 19.15 mA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
169 310 241 334
179 318 243 334
8 7.953 mA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
382 368 454 392
392 376 456 392
8 55.37 mW
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
381 351 453 375
391 359 455 375
8 11.19 mA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
497 340 569 364
507 348 571 364
8 41.71 mA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
498 355 554 379
508 363 556 379
6 501 mW
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
635 150 707 174
645 158 709 174
8 26.67 mA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
633 168 689 192
643 176 691 192
6 640 mW
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
384 335 448 359
394 343 450 359
7 4.947 V
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
497 325 561 349
507 333 563 349
7 12.01 V
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
635 130 675 154
645 138 677 154
4 24 V
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
4523550 1210432 100 100 0 0
0 0 0 0
11 120 172 190
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12401 0
4 2 5
1
255 87
0 5 0 0 2	3 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
