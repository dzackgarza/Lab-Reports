CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
40 0 30 150 9
36 70 1280 984
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
36 70 1280 984
144179218 0
0
6 Title:
5 Name:
0
0
0
12
11 Multimeter~
205 163 314 0 21 21
0 3 5 6 2 0 0 0 0 0
32 50 46 57 57 57 32 86 0 0
0 82
0
0 0 16464 180
8 100.0Meg
-29 -19 27 -11
3 MM0
-12 -29 9 -21
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
1 R
8953 0 0
0
0
7 Ground~
168 55 307 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4441 0 0
0
0
9 V Source~
197 56 220 0 2 5
0 4 2
0
0 0 17264 0
2 5V
16 0 30 8
3 Vs1
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
3618 0 0
0
0
13 Var Resistor~
219 169 228 0 3 7
0 4 3 2
0
0 0 848 270
8 100k 40%
-64 -4 -8 4
2 R1
-43 -14 -29 -6
0
0
32 %DA %1 %2 40000
%DB %2 %3 60000
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
82 0 0 0 1 0 0 0
1 R
6153 0 0
0
0
7 ADC0800
219 327 220 0 18 37
0 7 8 9 10 11 12 13 14 15
16 17 3 18 19 20 21 22 23
0
0 0 13008 0
7 ADC0800
-25 -56 24 -48
2 U1
-7 -56 7 -48
0
0
68 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %10 %11 %12 %13 %14 %15 %16 %17 %18 %S
0
0
5 DIP18
37

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 1
2 3 4 5 6 7 8 9 10 11
12 13 14 15 16 17 18 0
88 0 0 512 1 0 0 0
1 U
5394 0 0
0
0
4 LED~
171 1062 372 0 1 2
10 24
0
0 0 880 0
4 LED1
17 0 45 8
2 D7
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 512 0 0 0 0
1 D
7734 0 0
0
0
4 LED~
171 992 372 0 1 2
10 25
0
0 0 880 0
4 LED1
17 0 45 8
2 D6
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 512 0 0 0 0
1 D
9914 0 0
0
0
4 LED~
171 921 370 0 1 2
10 26
0
0 0 880 0
4 LED1
17 0 45 8
2 D5
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 512 0 0 0 0
1 D
3747 0 0
0
0
4 LED~
171 847 367 0 1 2
10 27
0
0 0 880 0
4 LED1
17 0 45 8
2 D4
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 512 0 0 0 0
1 D
3549 0 0
0
0
4 LED~
171 775 365 0 1 2
10 28
0
0 0 880 0
4 LED1
17 0 45 8
2 D3
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 512 0 0 0 0
1 D
7931 0 0
0
0
4 LED~
171 697 366 0 1 2
10 29
0
0 0 880 0
4 LED1
17 0 45 8
2 D2
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 512 0 0 0 0
1 D
9325 0 0
0
0
4 LED~
171 608 362 0 1 2
10 30
0
0 0 880 0
4 LED1
17 0 45 8
2 D1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 512 0 0 0 0
1 D
8903 0 0
0
0
6
4 0 2 0 0 4096 0 1 0 0 5 2
136 305
136 272
1 0 3 0 0 4096 0 1 0 0 3 2
186 305
231 305
2 12 3 0 0 12416 0 4 5 0 0 6
177 222
231 222
231 305
398 305
398 247
360 247
1 1 4 0 0 8320 0 4 3 0 0 4
165 206
165 173
56 173
56 199
3 0 2 0 0 8320 0 4 0 0 6 3
165 242
165 272
55 272
2 1 2 0 0 0 0 3 2 0 0 3
56 241
55 241
55 301
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
3015704 1079360 100 100 0 0
0 0 0 0
296 172 457 242
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12401 0
4 1 2
1
196 222
0 3 0 0 1	0 3 0 0
1704948 8550464 100 100 0 0
77 66 1247 366
-75 709 1205 1166
1247 66
77 66
1247 66
1247 366
0 0
5e-006 0 0.3 -0.3 5e-006 5e-006
12401 0
4 1e-006 2
1
154 272
0 2 0 0 2	0 5 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
