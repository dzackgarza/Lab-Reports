CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
180 0 30 100 9
112 110 1410 763
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
112 110 1410 763
144179218 0
0
6 Title:
5 Name:
0
0
0
8
9 Resistor~
219 230 149 0 1 5
0 0
0
0 0 864 0
3 10k
-10 -14 11 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8953 0 0
0
0
10 Capacitor~
219 163 148 0 1 5
0 0
0
0 0 832 0
5 150pF
-18 -18 17 -10
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
4441 0 0
0
0
7 Ground~
168 57 241 0 1 3
0 0
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3618 0 0
0
0
9 V Source~
197 149 395 0 1 5
0 0
0
0 0 17248 0
2 5V
17 0 31 8
3 Vs1
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
6153 0 0
0
0
13 Var Resistor~
219 192 280 0 1 7
0 0
0
0 0 832 0
7 10k 40%
-25 18 24 26
2 R1
-7 8 7 16
0
0
26 %DA %1 %2 4K
%DB %2 %3 6K
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
82 0 0 0 0 0 0 0
1 R
5394 0 0
0
0
7 Ground~
168 298 491 0 1 3
0 0
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7734 0 0
0
0
13 Logic Switch~
5 387 198 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
9914 0 0
0
0
7 ADC0800
219 608 223 0 1 37
0 0
0
0 0 12992 0
7 ADC0800
-25 -56 24 -48
2 U2
-7 -56 7 -48
0
0
68 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %10 %11 %12 %13 %14 %15 %16 %17 %18 %S
0
0
5 DIP18
37

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 1
2 3 4 5 6 7 8 9 10 11
12 13 14 15 16 17 18 0
88 0 0 0 1 0 0 0
1 U
3747 0 0
0
0
16
7 0 0 0 0 0 0 8 0 0 4 3
575 250
378 250
378 338
6 9 0 0 0 0 0 8 8 0 0 4
575 241
547 241
547 268
575 268
10 0 0 0 0 0 0 8 0 0 4 3
641 268
654 268
654 338
0 12 0 0 0 0 0 0 8 6 0 4
149 338
713 338
713 250
641 250
3 15 0 0 0 0 0 5 8 0 0 6
210 280
263 280
263 398
727 398
727 223
641 223
1 1 0 0 0 0 0 4 5 0 0 3
149 374
149 280
174 280
1 2 0 0 0 0 0 6 4 0 0 3
298 485
149 485
149 416
5 0 0 0 0 0 0 8 0 0 16 3
575 232
352 232
352 485
4 0 0 0 0 0 0 8 0 0 16 5
575 223
451 223
451 146
835 146
835 485
3 0 0 0 0 0 0 8 0 0 16 5
575 214
474 214
474 127
860 127
860 485
2 0 0 0 0 0 0 8 0 0 16 5
575 205
494 205
494 116
883 116
883 485
1 0 0 0 0 0 0 8 0 0 16 5
575 196
514 196
514 104
904 104
904 485
17 0 0 0 0 0 0 8 0 0 16 3
641 205
926 205
926 485
16 0 0 0 0 0 0 8 0 0 16 3
641 214
946 214
946 485
14 0 0 0 0 0 0 8 0 0 16 3
641 232
967 232
967 485
1 13 0 0 0 0 0 6 8 0 0 4
298 485
985 485
985 241
641 241
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
