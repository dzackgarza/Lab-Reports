CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
80 140 30 200 9
0 67 1280 411
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 67 1280 411
144179218 256
0
6 Title:
5 Name:
0
0
0
5
7 Ground~
168 324 315 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8953 0 0
0
0
9 Inductor~
219 468 225 0 2 5
0 4 3
0
0 0 848 270
4 17mH
9 -4 37 4
2 L1
10 -14 24 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
4441 0 0
0
0
10 Capacitor~
219 387 279 0 2 5
0 3 2
0
0 0 848 180
5 220uF
-18 -18 17 -10
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3618 0 0
0
0
11 Signal Gen~
195 288 225 0 19 64
0 5 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1203982336 0 1086324736
20
1 100000 0 6 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
5 -6/6V
-18 -30 17 -22
2 Vs
-7 -40 7 -32
0
0
38 %D %1 %2 DC 0 SIN(0 6 100k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
6153 0 0
0
0
9 Resistor~
219 387 171 0 2 5
0 5 4
0
0 0 880 0
3 12k
-10 -14 11 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5394 0 0
0
0
5
1 0 2 0 0 4096 0 1 0 0 2 2
324 309
324 279
2 2 2 0 0 4224 0 3 4 0 0 3
378 279
319 279
319 230
2 1 3 0 0 8320 0 2 3 0 0 3
468 243
468 279
396 279
2 1 4 0 0 4224 0 5 2 0 0 3
405 171
468 171
468 207
1 1 5 0 0 8320 0 4 5 0 0 3
319 220
319 171
369 171
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-005 2e-007 2e-007
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
459140 1210432 100 100 0 0
0 0 0 0
0 67 138 122
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12401 0
4 1 0.1
1
345 279
0 2 0 0 1	0 2 0 0
393602 276986432 100 100 0 0
66 61 1236 271
0 411 1280 755
1236 61
66 61
1236 61
1236 271
0 0
5e-005 0 5e-005 0 5e-005 5e-005
12409 0
4 1e-005 3
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
