CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
20 140 30 100 9
0 71 1366 768
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1366 768
177209362 0
0
6 Title:
5 Name:
0
0
0
40
4 LED~
171 1193 552 0 2 2
10 12 3
0
0 0 880 0
4 LED1
17 0 45 8
2 D9
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
8953 0 0
0
0
4 LED~
171 1154 555 0 2 2
10 10 3
0
0 0 880 0
4 LED1
17 0 45 8
2 D8
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
4441 0 0
0
0
4 LED~
171 1111 555 0 2 2
10 9 3
0
0 0 880 0
4 LED1
17 0 45 8
2 D7
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
3618 0 0
0
0
4 LED~
171 1071 556 0 2 2
10 8 3
0
0 0 880 0
4 LED1
17 0 45 8
2 D6
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
6153 0 0
0
0
4 LED~
171 1032 556 0 2 2
10 11 3
0
0 0 880 0
4 LED1
17 0 45 8
2 D5
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
5394 0 0
0
0
4 LED~
171 994 555 0 2 2
10 7 3
0
0 0 880 0
4 LED1
17 0 45 8
2 D4
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
7734 0 0
0
0
4 LED~
171 961 554 0 2 2
10 6 3
0
0 0 880 0
4 LED1
17 0 45 8
2 D3
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
9914 0 0
0
0
4 LED~
171 924 554 0 2 2
10 5 3
0
0 0 880 0
4 LED1
17 0 45 8
2 D2
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
3747 0 0
0
0
4 LED~
171 867 559 0 2 2
10 29 3
0
0 0 880 0
4 LED1
17 0 45 8
2 D1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
3549 0 0
0
0
7 Ground~
168 145 354 0 1 3
0 31
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7931 0 0
0
0
6 74LS83
105 808 177 0 14 29
0 31 31 31 31 19 18 17 16 31
8 9 10 12 30
0
0 0 13040 0
7 74LS83A
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
9325 0 0
0
0
6 74LS83
105 816 452 0 14 29
0 31 31 31 31 27 26 25 24 30
5 6 7 11 29
0
0 0 13040 0
7 74LS83A
-24 -60 25 -52
2 U3
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
8903 0 0
0
0
12 SPDT Switch~
164 288 344 0 3 11
0 31 39 31
0
0 0 5488 0
3 ADD
-11 12 10 20
2 SS
-7 -25 7 -17
8 SUBTRACT
-25 -19 31 -11
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 -1 0
1 S
3834 0 0
0
0
9 2-In XOR~
219 501 214 0 3 22
0 31 31 27
0
0 0 624 0
4 4070
-14 -24 14 -16
3 U4D
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 4 2 0
1 U
3363 0 0
0
0
9 2-In XOR~
219 499 268 0 3 22
0 31 31 26
0
0 0 624 0
4 4070
-14 -24 14 -16
3 U4C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 3 2 0
1 U
7668 0 0
0
0
9 2-In XOR~
219 503 319 0 3 22
0 31 31 25
0
0 0 624 0
4 4070
-14 -24 14 -16
3 U4B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 2 2 0
1 U
4718 0 0
0
0
9 2-In XOR~
219 503 399 0 3 22
0 31 31 24
0
0 0 624 0
4 4070
-14 -24 14 -16
3 U4A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 1 2 0
1 U
3874 0 0
0
0
9 2-In XOR~
219 503 455 0 3 22
0 31 31 19
0
0 0 624 0
4 4070
-14 -24 14 -16
3 U2D
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 4 1 0
1 U
6671 0 0
0
0
9 2-In XOR~
219 504 521 0 3 22
0 31 31 18
0
0 0 624 0
4 4070
-14 -24 14 -16
3 U2C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 3 1 0
1 U
3789 0 0
0
0
9 2-In XOR~
219 507 586 0 3 22
0 31 31 17
0
0 0 624 0
4 4070
-14 -24 14 -16
3 U2B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 2 1 0
1 U
4871 0 0
0
0
9 V Source~
197 68 630 0 2 5
0 39 31
0
0 0 17264 0
3 10V
13 0 34 8
3 Vs1
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
3750 0 0
0
0
12 SPDT Switch~
164 179 296 0 3 11
0 31 39 31
0
0 0 4720 0
0
2 A1
-8 -15 6 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
8778 0 0
0
0
12 SPDT Switch~
164 180 267 0 3 11
0 31 39 31
0
0 0 4720 0
0
2 A2
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
538 0 0
0
0
12 SPDT Switch~
164 187 242 0 3 11
0 31 39 31
0
0 0 4720 0
0
2 A3
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
6843 0 0
0
0
12 SPDT Switch~
164 187 213 0 3 11
0 31 39 31
0
0 0 4720 0
0
2 A4
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
3136 0 0
0
0
12 SPDT Switch~
164 182 183 0 3 11
0 31 39 31
0
0 0 4720 0
0
2 A5
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
5950 0 0
0
0
12 SPDT Switch~
164 185 156 0 3 11
0 31 39 31
0
0 0 4720 0
0
2 A6
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
5670 0 0
0
0
12 SPDT Switch~
164 186 125 0 3 11
0 31 39 31
0
0 0 4720 0
0
2 A7
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
6828 0 0
0
0
12 SPDT Switch~
164 184 95 0 3 11
0 31 39 31
0
0 0 4720 0
0
2 A8
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
6735 0 0
0
0
12 SPDT Switch~
164 185 558 0 3 11
0 31 39 31
0
0 0 4720 0
0
2 B2
-8 -16 6 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
8365 0 0
0
0
12 SPDT Switch~
164 184 529 0 3 11
0 31 39 31
0
0 0 4720 0
0
2 B3
-8 -16 6 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
4132 0 0
0
0
12 SPDT Switch~
164 183 503 0 3 11
0 31 39 31
0
0 0 4720 0
0
2 B4
-8 -16 6 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
4551 0 0
0
0
12 SPDT Switch~
164 183 476 0 3 11
0 31 39 31
0
0 0 4720 0
0
2 B5
-8 -16 6 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
3635 0 0
0
0
12 SPDT Switch~
164 181 447 0 3 11
0 31 39 31
0
0 0 4720 0
0
2 B6
-8 -16 6 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
3973 0 0
0
0
12 SPDT Switch~
164 183 419 0 3 11
0 31 39 31
0
0 0 4720 0
0
2 B7
-8 -16 6 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
3851 0 0
0
0
12 SPDT Switch~
164 182 391 0 3 11
0 31 39 31
0
0 0 4720 0
0
2 B8
-8 -16 6 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
8383 0 0
0
0
12 SPDT Switch~
164 184 591 0 3 11
0 31 39 31
0
0 0 4720 0
0
2 B1
-8 -16 6 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
9334 0 0
0
0
9 2-In XOR~
219 506 639 0 3 22
0 31 31 16
0
0 0 624 0
4 4070
-14 -24 14 -16
3 U2A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 1096765229
65 0 0 0 4 1 1 0
1 U
7471 0 0
0
0
7 Ground~
168 120 670 0 1 3
0 31
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3334 0 0
0
0
9 Resistor~
219 781 664 0 3 5
0 31 3 -1
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3559 0 0
0
0
90
2 2 3 0 0 4224 0 40 1 0 0 3
799 664
1193 664
1193 562
2 0 3 0 0 0 0 9 0 0 1 2
867 569
867 664
2 0 3 0 0 0 0 8 0 0 1 2
924 564
924 664
2 0 3 0 0 0 0 7 0 0 1 2
961 564
961 664
2 0 3 0 0 0 0 6 0 0 1 2
994 565
994 664
2 0 3 0 0 0 0 5 0 0 1 2
1032 566
1032 664
2 0 3 0 0 0 0 4 0 0 1 2
1071 566
1071 664
2 0 3 0 0 0 0 3 0 0 1 2
1111 565
1111 664
2 0 3 0 0 0 0 2 0 0 1 2
1154 565
1154 664
1 1 31 0 0 4224 4 29 12 0 0 4
201 95
741 95
741 416
784 416
1 0 31 0 0 0 2 10 0 0 48 2
145 348
145 348
1 1 31 0 0 4224 2 0 40 58 0 2
120 664
763 664
10 1 5 0 0 8320 0 12 8 0 0 3
848 443
924 443
924 544
11 1 6 0 0 4224 0 12 7 0 0 3
848 452
961 452
961 544
12 1 7 0 0 4224 0 12 6 0 0 4
848 461
995 461
995 545
994 545
10 1 8 0 0 8320 0 11 4 0 0 3
840 168
1071 168
1071 546
11 1 9 0 0 8320 0 11 3 0 0 3
840 177
1111 177
1111 545
12 1 10 0 0 8320 0 11 2 0 0 3
840 186
1154 186
1154 545
13 1 11 0 0 4224 0 12 5 0 0 3
848 470
1032 470
1032 546
13 1 12 0 0 4224 0 11 1 0 0 3
840 195
1193 195
1193 542
3 0 31 0 0 0 2 34 0 0 58 2
164 451
125 451
2 1 31 0 0 12416 13 12 28 0 0 6
784 425
725 425
725 107
221 107
221 125
203 125
3 1 31 0 0 12416 14 12 27 0 0 6
784 434
711 434
711 120
236 120
236 156
202 156
4 1 31 0 0 12416 15 12 26 0 0 6
784 443
699 443
699 131
249 131
249 183
199 183
3 8 16 0 0 8320 0 38 11 0 0 4
539 639
644 639
644 204
776 204
7 3 17 0 0 8320 0 11 20 0 0 4
776 195
631 195
631 586
540 586
3 6 18 0 0 8320 0 19 11 0 0 4
537 521
618 521
618 186
776 186
5 3 19 0 0 8320 0 11 18 0 0 6
776 177
606 177
606 439
547 439
547 455
536 455
1 1 31 0 0 4224 20 11 25 0 0 4
776 141
262 141
262 213
204 213
2 1 31 0 0 4224 21 11 24 0 0 4
776 150
286 150
286 242
204 242
3 1 31 0 0 4224 22 11 23 0 0 4
776 159
311 159
311 267
197 267
4 1 31 0 0 4224 23 11 22 0 0 4
776 168
331 168
331 296
196 296
8 3 24 0 0 4224 0 12 17 0 0 4
784 479
560 479
560 399
536 399
7 3 25 0 0 4224 0 12 16 0 0 4
784 470
572 470
572 319
536 319
6 3 26 0 0 4224 0 12 15 0 0 4
784 461
583 461
583 268
532 268
5 3 27 0 0 8320 0 12 14 0 0 4
784 452
593 452
593 214
534 214
0 9 31 0 0 4224 28 0 11 54 0 4
437 344
686 344
686 222
776 222
14 1 29 0 0 8320 0 12 9 0 0 3
848 497
867 497
867 549
14 9 30 0 0 12416 0 11 12 0 0 6
840 222
852 222
852 377
685 377
685 497
784 497
2 1 31 0 0 12416 0 38 37 0 0 4
490 648
400 648
400 591
201 591
2 1 31 0 0 12416 32 20 30 0 0 4
491 595
416 595
416 558
202 558
2 1 31 0 0 8320 33 19 31 0 0 3
488 530
488 529
201 529
2 1 31 0 0 12416 34 18 32 0 0 4
487 464
415 464
415 503
200 503
2 1 31 0 0 12416 35 17 33 0 0 4
487 408
397 408
397 476
200 476
2 1 31 0 0 12416 36 16 34 0 0 4
487 328
380 328
380 447
198 447
2 1 31 0 0 12416 37 15 35 0 0 4
483 277
364 277
364 419
200 419
1 2 31 0 0 8320 38 36 14 0 0 4
199 391
351 391
351 223
485 223
3 0 31 0 0 0 2 13 0 0 83 2
271 348
125 348
0 2 39 0 0 4096 0 0 13 72 0 3
68 339
271 339
271 340
0 1 31 0 0 0 28 0 38 51 0 3
437 577
437 630
490 630
1 0 31 0 0 0 28 20 0 0 52 3
491 577
437 577
437 512
1 0 31 0 0 0 28 19 0 0 53 3
488 512
437 512
437 446
1 0 31 0 0 0 28 18 0 0 54 3
487 446
437 446
437 390
1 0 31 0 0 0 28 17 0 0 57 3
487 390
437 390
437 344
1 0 31 0 0 0 28 16 0 0 57 2
487 310
437 310
1 0 31 0 0 0 28 15 0 0 57 2
483 259
437 259
1 1 31 0 0 0 28 14 13 0 0 4
485 205
437 205
437 344
305 344
0 1 31 0 0 0 2 0 39 0 0 3
125 375
125 664
120 664
3 0 31 0 0 0 2 37 0 0 58 2
167 595
125 595
3 0 31 0 0 0 2 30 0 0 58 2
168 562
125 562
3 0 31 0 0 0 2 31 0 0 58 2
167 533
125 533
3 0 31 0 0 0 2 32 0 0 58 2
166 507
125 507
3 0 31 0 0 0 2 33 0 0 58 2
166 480
125 480
3 0 31 0 0 0 2 35 0 0 58 2
166 423
125 423
3 0 31 0 0 0 2 36 0 0 58 2
165 395
125 395
2 0 39 0 0 0 0 36 0 0 72 2
165 387
68 387
2 0 39 0 0 0 0 35 0 0 72 2
166 415
68 415
2 0 39 0 0 0 0 34 0 0 72 2
164 443
68 443
2 0 39 0 0 0 0 33 0 0 72 2
166 472
68 472
2 0 39 0 0 0 0 32 0 0 72 2
166 499
68 499
2 0 39 0 0 0 0 31 0 0 72 2
167 525
68 525
2 2 39 0 0 8320 0 30 29 0 0 4
168 554
68 554
68 91
167 91
2 0 39 0 0 0 0 37 0 0 75 2
167 587
68 587
1 2 31 0 0 0 2 39 21 0 0 3
120 664
68 664
68 651
1 0 39 0 0 0 0 21 0 0 72 3
68 609
68 554
69 554
3 0 31 0 0 0 2 22 0 0 83 2
162 300
125 300
3 0 31 0 0 0 2 23 0 0 83 2
163 271
125 271
3 0 31 0 0 0 2 24 0 0 83 2
170 246
125 246
3 0 31 0 0 0 2 25 0 0 83 2
170 217
125 217
3 0 31 0 0 0 2 26 0 0 83 2
165 187
125 187
3 0 31 0 0 0 2 27 0 0 83 2
168 160
125 160
3 0 31 0 0 0 2 28 0 0 83 2
169 129
125 129
3 0 31 0 0 0 2 29 0 0 0 3
167 99
125 99
125 376
2 0 39 0 0 0 0 22 0 0 72 2
162 292
68 292
2 0 39 0 0 0 0 23 0 0 72 2
163 263
68 263
2 0 39 0 0 0 0 24 0 0 72 2
170 238
68 238
2 0 39 0 0 0 0 25 0 0 72 2
170 209
68 209
2 0 39 0 0 0 0 26 0 0 72 2
165 179
68 179
2 0 39 0 0 0 0 27 0 0 72 2
168 152
68 152
2 0 39 0 0 0 0 28 0 0 72 2
169 121
68 121
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
1312660 1210432 100 100 0 0
0 0 0 0
1 66 162 136
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12401 0
4 2 2
1
791 284
0 11 0 0 2	0 91 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
