CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 370 30 100 9
0 70 1275 793
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 70 1275 793
177209362 0
0
6 Title:
5 Name:
0
0
0
48
7 Ground~
168 262 996 0 1 3
0 53
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8953 0 0
0
0
9 V Source~
197 264 946 0 2 5
0 3 53
0
0 0 17264 0
3 -5V
13 0 34 8
3 Vs2
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
4441 0 0
0
0
7 Ground~
168 609 749 0 1 3
0 53
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3618 0 0
0
0
10 Capacitor~
219 514 879 0 2 5
0 53 6
0
0 0 848 90
5 150uF
4 0 39 8
2 C1
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6153 0 0
0
0
7 ADC0800
219 317 742 0 18 37
0 12 11 10 9 53 5 54 3 5
54 7 8 16 15 54 14 13 53
0
0 0 13008 0
7 ADC0800
-25 -56 24 -48
2 U5
-7 -56 7 -48
0
0
68 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %10 %11 %12 %13 %14 %15 %16 %17 %18 %S
0
0
5 DIP18
37

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 1
2 3 4 5 6 7 8 9 10 11
12 13 14 15 16 17 18 0
88 0 0 0 1 0 0 0
1 U
5394 0 0
0
0
13 Var Resistor~
219 73 817 0 3 7
0 54 8 53
0
0 0 848 270
6 1k 10%
-58 -4 -16 4
2 R2
-43 -14 -29 -6
0
0
28 %DA %1 %2 100
%DB %2 %3 900
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
82 0 0 0 1 0 0 0
1 R
7734 0 0
0
0
11 Multimeter~
205 122 962 0 21 21
0 8 45 46 53 0 0 0 0 0
78 79 32 68 65 84 65 32 0 0
0 82
0
0 0 16464 180
8 100.0Meg
-29 -19 27 -11
3 MM0
-12 -29 9 -21
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
1 R
9914 0 0
0
0
4 LED~
171 1072 560 0 2 2
10 22 18
0
0 0 864 0
4 LED1
17 0 45 8
2 D9
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3747 0 0
0
0
4 LED~
171 1112 625 0 2 2
10 23 18
0
0 0 864 0
4 LED1
17 0 45 8
2 D8
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3549 0 0
0
0
4 LED~
171 1151 626 0 2 2
10 24 18
0
0 0 864 0
4 LED1
17 0 45 8
2 D7
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
7931 0 0
0
0
4 LED~
171 1191 627 0 2 2
10 26 18
0
0 0 864 0
4 LED1
17 0 45 8
2 D6
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
9325 0 0
0
0
4 LED~
171 1032 620 0 2 2
10 25 18
0
0 0 864 0
4 LED1
17 0 45 8
2 D5
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
8903 0 0
0
0
4 LED~
171 997 578 0 2 2
10 19 18
0
0 0 864 0
4 LED1
17 0 45 8
2 D4
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3834 0 0
0
0
4 LED~
171 960 573 0 2 2
10 17 18
0
0 0 864 0
4 LED1
17 0 45 8
2 D3
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3363 0 0
0
0
4 LED~
171 920 595 0 2 2
10 20 18
0
0 0 864 0
4 LED1
17 0 45 8
2 D2
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
7668 0 0
0
0
4 LED~
171 873 591 0 2 2
10 21 18
0
0 0 864 0
4 LED1
17 0 45 8
2 D1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
4718 0 0
0
0
7 Ground~
168 145 354 0 1 3
0 53
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3874 0 0
0
0
6 74LS83
105 808 177 0 14 29
0 53 53 53 53 34 33 32 31 53
22 23 24 26 44
0
0 0 13040 0
7 74LS83A
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
6671 0 0
0
0
6 74LS83
105 813 301 0 14 29
0 53 53 53 53 42 41 40 39 44
20 17 19 25 21
0
0 0 13040 0
7 74LS83A
-24 -60 25 -52
2 U3
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
3789 0 0
0
0
12 SPDT Switch~
164 288 344 0 3 11
0 53 54 53
0
0 0 5488 0
3 ADD
-11 12 10 20
2 SS
-7 -25 7 -17
8 SUBTRACT
-25 -19 31 -11
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 -1 0
1 S
4871 0 0
0
0
9 2-In XOR~
219 501 214 0 3 22
0 53 9 42
0
0 0 624 0
4 4070
-14 -24 14 -16
3 U4D
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 4 2 0
1 U
3750 0 0
0
0
9 2-In XOR~
219 499 268 0 3 22
0 53 10 41
0
0 0 624 0
4 4070
-14 -24 14 -16
3 U4C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 3 2 0
1 U
8778 0 0
0
0
9 2-In XOR~
219 503 319 0 3 22
0 53 11 40
0
0 0 624 0
4 4070
-14 -24 14 -16
3 U4B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 2 2 0
1 U
538 0 0
0
0
9 2-In XOR~
219 503 399 0 3 22
0 53 12 39
0
0 0 624 0
4 4070
-14 -24 14 -16
3 U4A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 1 2 0
1 U
6843 0 0
0
0
9 2-In XOR~
219 503 455 0 3 22
0 53 13 34
0
0 0 624 0
4 4070
-14 -24 14 -16
3 U2D
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 4 1 0
1 U
3136 0 0
0
0
9 2-In XOR~
219 504 521 0 3 22
0 53 14 33
0
0 0 624 0
4 4070
-14 -24 14 -16
3 U2C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 3 1 0
1 U
5950 0 0
0
0
9 2-In XOR~
219 507 586 0 3 22
0 53 15 32
0
0 0 624 0
4 4070
-14 -24 14 -16
3 U2B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 2 1 0
1 U
5670 0 0
0
0
9 V Source~
197 68 630 0 2 5
0 54 53
0
0 0 17264 0
2 5V
16 0 30 8
3 Vs1
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
6828 0 0
0
0
12 SPDT Switch~
164 179 296 0 3 11
0 53 54 53
0
0 0 4720 0
0
2 A1
-8 -15 6 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
6735 0 0
0
0
12 SPDT Switch~
164 180 267 0 3 11
0 53 54 53
0
0 0 4720 0
0
2 A2
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
8365 0 0
0
0
12 SPDT Switch~
164 187 242 0 3 11
0 53 54 53
0
0 0 4720 0
0
2 A3
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
4132 0 0
0
0
12 SPDT Switch~
164 187 213 0 3 11
0 53 54 53
0
0 0 4720 0
0
2 A4
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
4551 0 0
0
0
12 SPDT Switch~
164 182 183 0 3 11
0 53 54 53
0
0 0 4720 0
0
2 A5
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
3635 0 0
0
0
12 SPDT Switch~
164 185 156 0 3 11
0 53 54 53
0
0 0 4720 0
0
2 A6
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
3973 0 0
0
0
12 SPDT Switch~
164 186 125 0 3 11
0 53 54 53
0
0 0 4720 0
0
2 A7
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
3851 0 0
0
0
12 SPDT Switch~
164 184 95 0 3 11
0 53 54 53
0
0 0 4720 0
0
2 A8
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
8383 0 0
0
0
12 SPDT Switch~
164 185 558 0 10 11
0 47 54 53 0 0 0 0 0 0
1
0
0 0 4720 0
0
2 B2
-8 -16 6 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 512 1 0 0 0
1 S
9334 0 0
0
0
12 SPDT Switch~
164 184 529 0 10 11
0 48 54 53 0 0 0 0 0 0
1
0
0 0 4720 0
0
2 B3
-8 -16 6 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 512 1 0 0 0
1 S
7471 0 0
0
0
12 SPDT Switch~
164 183 503 0 10 11
0 49 54 53 0 0 0 0 0 0
1
0
0 0 4720 0
0
2 B4
-8 -16 6 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 512 1 0 0 0
1 S
3334 0 0
0
0
12 SPDT Switch~
164 183 476 0 10 11
0 50 54 53 0 0 0 0 0 0
1
0
0 0 4720 0
0
2 B5
-8 -16 6 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 512 1 0 0 0
1 S
3559 0 0
0
0
12 SPDT Switch~
164 181 447 0 10 11
0 51 54 53 0 0 0 0 0 0
1
0
0 0 4720 0
0
2 B6
-8 -16 6 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 512 1 0 0 0
1 S
984 0 0
0
0
12 SPDT Switch~
164 183 419 0 3 11
0 52 54 53
0
0 0 4720 0
0
2 B7
-8 -16 6 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 512 1 0 0 0
1 S
7557 0 0
0
0
12 SPDT Switch~
164 182 391 0 3 11
0 53 54 53
0
0 0 4720 0
0
2 B8
-8 -16 6 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 512 1 0 0 0
1 S
3146 0 0
0
0
12 SPDT Switch~
164 184 591 0 10 11
0 54 54 53 0 0 0 0 0 0
1
0
0 0 4720 0
0
2 B1
-8 -16 6 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 512 1 0 0 0
1 S
5687 0 0
0
0
9 2-In XOR~
219 506 639 0 3 22
0 53 16 31
0
0 0 624 0
4 4070
-14 -24 14 -16
3 U2A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 1096765229
65 0 0 0 4 1 1 0
1 U
7939 0 0
0
0
7 Ground~
168 126 756 0 1 3
0 53
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3308 0 0
0
0
9 Resistor~
219 514 829 0 2 5
0 6 7
0
0 0 880 90
3 10k
5 0 26 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3408 0 0
0
0
9 Resistor~
219 925 684 0 3 5
0 53 18 -1
0
0 0 880 0
3 300
-10 -14 11 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9773 0 0
0
0
114
2 1 53 0 0 8192 2 2 1 0 0 3
264 967
262 967
262 990
1 8 3 0 0 4224 0 2 5 0 0 3
264 925
264 778
284 778
0 5 53 0 0 4096 2 0 5 83 0 4
126 740
218 740
218 751
284 751
15 0 54 0 0 4096 4 5 0 0 8 4
350 742
464 742
464 846
385 846
18 1 53 0 0 4096 2 5 3 0 0 3
350 715
609 715
609 743
9 6 5 0 0 8320 0 5 5 0 0 4
284 787
260 787
260 760
284 760
0 7 54 0 0 0 4 0 5 8 0 3
241 768
241 769
284 769
0 10 54 0 0 4112 4 0 5 16 0 6
29 768
241 768
241 852
385 852
385 787
350 787
1 0 53 0 0 4096 2 4 0 0 83 4
514 888
201 888
201 700
125 700
1 2 6 0 0 4224 0 47 4 0 0 2
514 847
514 870
11 2 7 0 0 4224 0 5 47 0 0 3
350 778
514 778
514 811
1 0 8 0 0 8192 0 7 0 0 14 3
145 953
164 953
164 811
4 0 53 0 0 0 2 7 0 0 15 3
95 953
69 953
69 897
2 12 8 0 0 4224 0 6 5 0 0 4
81 811
440 811
440 769
350 769
3 0 53 0 0 0 2 6 0 0 17 4
69 831
69 899
109 899
109 717
0 1 54 0 0 0 4 0 6 99 0 4
68 596
29 596
29 795
69 795
2 0 53 0 0 0 2 28 0 0 83 3
68 651
68 717
125 717
2 4 9 0 0 8320 0 21 5 0 0 6
485 223
350 223
350 553
237 553
237 742
284 742
2 3 10 0 0 8320 0 22 5 0 0 6
483 277
366 277
366 576
224 576
224 733
284 733
2 2 11 0 0 16512 0 23 5 0 0 6
487 328
396 328
396 469
265 469
265 724
284 724
2 1 12 0 0 8320 0 24 5 0 0 4
487 408
277 408
277 715
284 715
2 17 13 0 0 8320 0 25 5 0 0 4
487 464
408 464
408 724
350 724
2 16 14 0 0 8320 0 26 5 0 0 4
488 530
372 530
372 733
350 733
2 14 15 0 0 8320 0 27 5 0 0 4
491 595
356 595
356 751
350 751
2 13 16 0 0 8320 0 45 5 0 0 4
490 648
380 648
380 760
350 760
1 0 17 0 0 4096 0 14 0 0 48 2
960 563
960 571
0 0 18 0 0 4096 0 0 0 39 36 2
1062 673
1072 673
0 0 18 0 0 0 0 0 0 38 39 2
1053 666
1062 666
0 0 18 0 0 0 0 0 0 37 38 2
1044 675
1053 675
0 0 18 0 0 0 0 0 0 41 37 2
1035 667
1044 667
0 0 18 0 0 0 0 0 0 46 41 2
1026 674
1035 674
0 0 18 0 0 0 0 0 0 45 46 2
1017 666
1026 666
0 0 18 0 0 0 0 0 0 45 45 2
1008 676
1017 676
0 0 18 0 0 0 0 0 0 35 45 2
999 671
1008 671
2 2 18 0 0 16384 0 48 16 0 0 6
943 684
943 685
999 685
999 655
873 655
873 601
2 0 18 0 0 0 0 8 0 0 39 3
1072 570
1072 684
1062 684
2 0 18 0 0 0 0 9 0 0 41 5
1112 635
1112 646
1044 646
1044 685
1035 685
2 0 18 0 0 0 0 10 0 0 37 5
1151 636
1151 651
1053 651
1053 685
1044 685
2 0 18 0 0 8320 0 11 0 0 38 5
1191 637
1191 655
1062 655
1062 685
1053 685
1 12 19 0 0 4224 0 13 19 0 0 3
997 568
997 310
845 310
0 2 18 0 0 0 0 0 12 46 0 5
1026 685
1035 685
1035 637
1032 637
1032 630
10 1 20 0 0 8320 0 19 15 0 0 3
845 292
920 292
920 585
14 1 21 0 0 8320 0 19 16 0 0 3
845 346
873 346
873 581
0 1 53 0 0 12416 2 0 48 83 0 5
125 664
182 664
182 685
907 685
907 684
2 2 18 0 0 0 0 14 15 0 0 8
960 583
960 636
1017 636
1017 685
1008 685
1008 643
920 643
920 605
2 0 18 0 0 0 0 13 0 0 0 5
997 588
997 629
1026 629
1026 685
1017 685
1 0 53 0 0 0 2 17 0 0 73 2
145 348
145 348
11 1 17 0 0 8320 0 19 14 0 0 5
845 301
960 301
960 571
960 571
960 563
10 1 22 0 0 8320 0 18 8 0 0 3
840 168
1072 168
1072 550
11 1 23 0 0 8320 0 18 9 0 0 4
840 177
1111 177
1111 615
1112 615
12 1 24 0 0 8320 0 18 10 0 0 3
840 186
1151 186
1151 616
13 1 25 0 0 8320 0 19 12 0 0 3
845 319
1032 319
1032 610
13 1 26 0 0 8320 0 18 11 0 0 4
840 195
1190 195
1190 617
1191 617
3 0 53 0 0 0 2 41 0 0 83 2
164 451
125 451
1 1 53 0 0 4224 27 36 19 0 0 4
201 95
741 95
741 265
781 265
2 1 53 0 0 12416 28 19 35 0 0 6
781 274
725 274
725 107
221 107
221 125
203 125
3 1 53 0 0 12416 29 19 34 0 0 6
781 283
711 283
711 120
236 120
236 156
202 156
4 1 53 0 0 12416 30 19 33 0 0 6
781 292
699 292
699 131
249 131
249 183
199 183
3 8 31 0 0 8320 0 45 18 0 0 4
539 639
644 639
644 204
776 204
7 3 32 0 0 8320 0 18 27 0 0 4
776 195
631 195
631 586
540 586
3 6 33 0 0 8320 0 26 18 0 0 4
537 521
618 521
618 186
776 186
5 3 34 0 0 8320 0 18 25 0 0 6
776 177
606 177
606 439
547 439
547 455
536 455
1 1 53 0 0 4224 35 18 32 0 0 4
776 141
262 141
262 213
204 213
2 1 53 0 0 4224 36 18 31 0 0 4
776 150
286 150
286 242
204 242
3 1 53 0 0 4224 37 18 30 0 0 4
776 159
311 159
311 267
197 267
4 1 53 0 0 4224 38 18 29 0 0 4
776 168
331 168
331 296
196 296
8 3 39 0 0 4224 0 19 24 0 0 4
781 328
560 328
560 399
536 399
7 3 40 0 0 4224 0 19 23 0 0 2
781 319
536 319
6 3 41 0 0 4224 0 19 22 0 0 4
781 310
583 310
583 268
532 268
5 3 42 0 0 4224 0 19 21 0 0 4
781 301
593 301
593 214
534 214
0 9 53 0 0 4224 43 0 18 79 0 4
437 344
686 344
686 222
776 222
14 9 44 0 0 12416 0 18 19 0 0 6
840 222
852 222
852 377
685 377
685 346
781 346
3 0 53 0 0 0 2 20 0 0 107 2
271 348
125 348
0 2 54 0 0 0 4 0 20 97 0 3
68 339
271 339
271 340
0 1 53 0 0 0 43 0 45 76 0 3
437 577
437 630
490 630
1 0 53 0 0 0 43 27 0 0 77 3
491 577
437 577
437 512
1 0 53 0 0 0 43 26 0 0 78 3
488 512
437 512
437 446
1 0 53 0 0 0 43 25 0 0 79 3
487 446
437 446
437 390
1 0 53 0 0 0 43 24 0 0 82 3
487 390
437 390
437 344
1 0 53 0 0 0 43 23 0 0 82 2
487 310
437 310
1 0 53 0 0 0 43 22 0 0 82 2
483 259
437 259
1 1 53 0 0 0 43 21 20 0 0 4
485 205
437 205
437 344
305 344
0 1 53 0 0 0 2 0 46 0 0 4
125 375
125 717
126 717
126 750
3 0 53 0 0 0 2 44 0 0 83 2
167 595
125 595
3 0 53 0 0 0 2 37 0 0 83 2
168 562
125 562
3 0 53 0 0 0 2 38 0 0 83 2
167 533
125 533
3 0 53 0 0 0 2 39 0 0 83 2
166 507
125 507
3 0 53 0 0 0 2 40 0 0 83 2
166 480
125 480
3 0 53 0 0 0 2 42 0 0 83 2
166 423
125 423
3 0 53 0 0 0 2 43 0 0 83 2
165 395
125 395
2 0 54 0 0 0 4 43 0 0 97 2
165 387
68 387
2 0 54 0 0 0 4 42 0 0 97 2
166 415
68 415
2 0 54 0 0 0 4 41 0 0 97 2
164 443
68 443
2 0 54 0 0 0 4 40 0 0 97 2
166 472
68 472
2 0 54 0 0 0 4 39 0 0 97 2
166 499
68 499
2 0 54 0 0 0 4 38 0 0 97 2
167 525
68 525
2 2 54 0 0 8320 4 37 36 0 0 4
168 554
68 554
68 91
167 91
2 0 54 0 0 0 4 44 0 0 99 2
167 587
68 587
1 0 54 0 0 0 4 28 0 0 97 3
68 609
68 554
69 554
3 0 53 0 0 0 2 29 0 0 107 2
162 300
125 300
3 0 53 0 0 0 2 30 0 0 107 2
163 271
125 271
3 0 53 0 0 0 2 31 0 0 107 2
170 246
125 246
3 0 53 0 0 0 2 32 0 0 107 2
170 217
125 217
3 0 53 0 0 0 2 33 0 0 107 2
165 187
125 187
3 0 53 0 0 0 2 34 0 0 107 2
168 160
125 160
3 0 53 0 0 0 2 35 0 0 107 2
169 129
125 129
3 0 53 0 0 0 2 36 0 0 0 3
167 99
125 99
125 376
2 0 54 0 0 0 4 29 0 0 97 2
162 292
68 292
2 0 54 0 0 0 4 30 0 0 97 2
163 263
68 263
2 0 54 0 0 0 4 31 0 0 97 2
170 238
68 238
2 0 54 0 0 0 4 32 0 0 97 2
170 209
68 209
2 0 54 0 0 0 4 33 0 0 97 2
165 179
68 179
2 0 54 0 0 0 4 34 0 0 97 2
168 152
68 152
2 0 54 0 0 0 4 35 0 0 97 2
169 121
68 121
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
6030214 1210432 100 100 0 0
0 0 0 0
0 70 161 140
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12401 0
4 1 2
0
4195326 8550464 100 100 0 0
77 66 1247 366
0 527 1280 984
1247 66
77 66
1247 66
1247 366
0 0
5e-006 0 5e-006 0 5e-006 5e-006
12385 0
4 1e-006 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
